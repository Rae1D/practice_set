`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/08/05 09:40:54
// Design Name: 
// Module Name: add_zizhen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module add_zizhen(
   input clk,


    input data_in_valid,
    input [15:0]data_in_L_1_I ,
    input [15:0]data_in_L_1_Q ,
    input [15:0]data_in_L_2_I ,
    input [15:0]data_in_L_2_Q ,
    input [15:0]data_in_L_3_I ,
    input [15:0]data_in_L_3_Q ,
    input [15:0]data_in_L_4_I ,
    input [15:0]data_in_L_4_Q ,
    input [15:0]data_in_L_5_I ,
    input [15:0]data_in_L_5_Q ,
    input [15:0]data_in_L_6_I ,
    input [15:0]data_in_L_6_Q ,
    input [15:0]data_in_L_7_I ,
    input [15:0]data_in_L_7_Q ,
    input [15:0]data_in_L_8_I ,
    input [15:0]data_in_L_8_Q ,
    input [15:0]data_in_L_9_I ,
    input [15:0]data_in_L_9_Q ,
    input [15:0]data_in_L_10_I,
    input [15:0]data_in_L_10_Q,
    input [15:0]data_in_L_11_I,
    input [15:0]data_in_L_11_Q,
    input [15:0]data_in_L_12_I,
    input [15:0]data_in_L_12_Q,
    input [15:0]data_in_L_13_I,
    input [15:0]data_in_L_13_Q,
    input [15:0]data_in_L_14_I,
    input [15:0]data_in_L_14_Q,
    input [15:0]data_in_L_15_I,
    input [15:0]data_in_L_15_Q,
    input [15:0]data_in_L_16_I,
    input [15:0]data_in_L_16_Q,
    input [15:0]data_in_L_17_I,
    input [15:0]data_in_L_17_Q,
    input [15:0]data_in_L_18_I,
    input [15:0]data_in_L_18_Q,
    input [15:0]data_in_L_19_I,
    input [15:0]data_in_L_19_Q,
    input [15:0]data_in_L_20_I,
    input [15:0]data_in_L_20_Q,
    input [15:0]data_in_L_21_I,
    input [15:0]data_in_L_21_Q,
    input [15:0]data_in_L_22_I,
    input [15:0]data_in_L_22_Q,
    input [15:0]data_in_L_23_I,
    input [15:0]data_in_L_23_Q,
    input [15:0]data_in_L_24_I,
    input [15:0]data_in_L_24_Q,
    input [15:0]data_in_L_25_I,
    input [15:0]data_in_L_25_Q,
    input [15:0]data_in_L_26_I,
    input [15:0]data_in_L_26_Q,
    input [15:0]data_in_L_27_I,
    input [15:0]data_in_L_27_Q,
    input [15:0]data_in_L_28_I,
    input [15:0]data_in_L_28_Q,
    input [15:0]data_in_L_29_I,
    input [15:0]data_in_L_29_Q,
    input [15:0]data_in_L_30_I,
    input [15:0]data_in_L_30_Q,
    input [15:0]data_in_L_31_I,
    input [15:0]data_in_L_31_Q,
    input [15:0]data_in_L_32_I,
    input [15:0]data_in_L_32_Q,
    input [15:0]data_in_L_33_I,
    input [15:0]data_in_L_33_Q,
    input [15:0]data_in_L_34_I,
    input [15:0]data_in_L_34_Q,
    input [15:0]data_in_L_35_I,
    input [15:0]data_in_L_35_Q,
    input [15:0]data_in_L_36_I,
    input [15:0]data_in_L_36_Q,
    input [15:0]data_in_L_37_I,
    input [15:0]data_in_L_37_Q,
    input [15:0]data_in_L_38_I,
    input [15:0]data_in_L_38_Q,
    input [15:0]data_in_L_39_I,
    input [15:0]data_in_L_39_Q,
    input [15:0]data_in_L_40_I,
    input [15:0]data_in_L_40_Q,
    input [15:0]data_in_L_41_I,
    input [15:0]data_in_L_41_Q,
    input [15:0]data_in_L_42_I,
    input [15:0]data_in_L_42_Q,
    input [15:0]data_in_L_43_I,
    input [15:0]data_in_L_43_Q,
    input [15:0]data_in_L_44_I,
    input [15:0]data_in_L_44_Q,
    input [15:0]data_in_L_45_I,
    input [15:0]data_in_L_45_Q,
    input [15:0]data_in_L_46_I,
    input [15:0]data_in_L_46_Q,
    input [15:0]data_in_L_47_I,
    input [15:0]data_in_L_47_Q,
    input [15:0]data_in_L_48_I,
    input [15:0]data_in_L_48_Q,
    input [15:0]data_in_L_49_I,
    input [15:0]data_in_L_49_Q,
    input [15:0]data_in_L_50_I,
    input [15:0]data_in_L_50_Q,
    input [15:0]data_in_L_51_I,
    input [15:0]data_in_L_51_Q,
    input [15:0]data_in_L_52_I,
    input [15:0]data_in_L_52_Q,
    input [15:0]data_in_L_53_I,
    input [15:0]data_in_L_53_Q,
    input [15:0]data_in_L_54_I,
    input [15:0]data_in_L_54_Q,
    input [15:0]data_in_L_55_I,
    input [15:0]data_in_L_55_Q,
    input [15:0]data_in_L_56_I,
    input [15:0]data_in_L_56_Q,
    input [15:0]data_in_L_57_I,
    input [15:0]data_in_L_57_Q,
    input [15:0]data_in_L_58_I,
    input [15:0]data_in_L_58_Q,
    input [15:0]data_in_L_59_I,
    input [15:0]data_in_L_59_Q,
    input [15:0]data_in_L_60_I,
    input [15:0]data_in_L_60_Q,
    input [15:0]data_in_L_61_I,
    input [15:0]data_in_L_61_Q,
    input [15:0]data_in_L_62_I,
    input [15:0]data_in_L_62_Q,
    input [15:0]data_in_L_63_I,
    input [15:0]data_in_L_63_Q,
    input [15:0]data_in_L_64_I,
    input [15:0]data_in_L_64_Q,
    input [15:0]data_in_L_65_I,
    input [15:0]data_in_L_65_Q,
    input [15:0]data_in_L_66_I,
    input [15:0]data_in_L_66_Q,
    input [15:0]data_in_L_67_I,
    input [15:0]data_in_L_67_Q,
    input [15:0]data_in_L_68_I,
    input [15:0]data_in_L_68_Q,
    input [15:0]data_in_L_69_I,
    input [15:0]data_in_L_69_Q,
    input [15:0]data_in_L_70_I,
    input [15:0]data_in_L_70_Q,
    
    input [15:0]data_in_R_1_I ,
    input [15:0]data_in_R_1_Q ,
    input [15:0]data_in_R_2_I ,
    input [15:0]data_in_R_2_Q ,
    input [15:0]data_in_R_3_I ,
    input [15:0]data_in_R_3_Q ,
    input [15:0]data_in_R_4_I ,
    input [15:0]data_in_R_4_Q ,
    input [15:0]data_in_R_5_I ,
    input [15:0]data_in_R_5_Q ,
    input [15:0]data_in_R_6_I ,
    input [15:0]data_in_R_6_Q ,
    input [15:0]data_in_R_7_I ,
    input [15:0]data_in_R_7_Q ,
    input [15:0]data_in_R_8_I ,
    input [15:0]data_in_R_8_Q ,
    input [15:0]data_in_R_9_I ,
    input [15:0]data_in_R_9_Q ,
    input [15:0]data_in_R_10_I,
    input [15:0]data_in_R_10_Q,
    input [15:0]data_in_R_11_I,
    input [15:0]data_in_R_11_Q,
    input [15:0]data_in_R_12_I,
    input [15:0]data_in_R_12_Q,
    input [15:0]data_in_R_13_I,
    input [15:0]data_in_R_13_Q,
    input [15:0]data_in_R_14_I,
    input [15:0]data_in_R_14_Q,
    input [15:0]data_in_R_15_I,
    input [15:0]data_in_R_15_Q,
    input [15:0]data_in_R_16_I,
    input [15:0]data_in_R_16_Q,
    input [15:0]data_in_R_17_I,
    input [15:0]data_in_R_17_Q,
    input [15:0]data_in_R_18_I,
    input [15:0]data_in_R_18_Q,
    input [15:0]data_in_R_19_I,
    input [15:0]data_in_R_19_Q,
    input [15:0]data_in_R_20_I,
    input [15:0]data_in_R_20_Q,
    input [15:0]data_in_R_21_I,
    input [15:0]data_in_R_21_Q,
    input [15:0]data_in_R_22_I,
    input [15:0]data_in_R_22_Q,
    input [15:0]data_in_R_23_I,
    input [15:0]data_in_R_23_Q,
    input [15:0]data_in_R_24_I,
    input [15:0]data_in_R_24_Q,
    input [15:0]data_in_R_25_I,
    input [15:0]data_in_R_25_Q,
    input [15:0]data_in_R_26_I,
    input [15:0]data_in_R_26_Q,
    input [15:0]data_in_R_27_I,
    input [15:0]data_in_R_27_Q,
    input [15:0]data_in_R_28_I,
    input [15:0]data_in_R_28_Q,
    input [15:0]data_in_R_29_I,
    input [15:0]data_in_R_29_Q,
    input [15:0]data_in_R_30_I,
    input [15:0]data_in_R_30_Q,
    input [15:0]data_in_R_31_I,
    input [15:0]data_in_R_31_Q,
    input [15:0]data_in_R_32_I,
    input [15:0]data_in_R_32_Q,
    input [15:0]data_in_R_33_I,
    input [15:0]data_in_R_33_Q,
    input [15:0]data_in_R_34_I,
    input [15:0]data_in_R_34_Q,
    input [15:0]data_in_R_35_I,
    input [15:0]data_in_R_35_Q,
    input [15:0]data_in_R_36_I,
    input [15:0]data_in_R_36_Q,
    input [15:0]data_in_R_37_I,
    input [15:0]data_in_R_37_Q,
    input [15:0]data_in_R_38_I,
    input [15:0]data_in_R_38_Q,
    input [15:0]data_in_R_39_I,
    input [15:0]data_in_R_39_Q,
    input [15:0]data_in_R_40_I,
    input [15:0]data_in_R_40_Q,
    input [15:0]data_in_R_41_I,
    input [15:0]data_in_R_41_Q,
    input [15:0]data_in_R_42_I,
    input [15:0]data_in_R_42_Q,
    input [15:0]data_in_R_43_I,
    input [15:0]data_in_R_43_Q,
    input [15:0]data_in_R_44_I,
    input [15:0]data_in_R_44_Q,
    input [15:0]data_in_R_45_I,
    input [15:0]data_in_R_45_Q,
    input [15:0]data_in_R_46_I,
    input [15:0]data_in_R_46_Q,
    input [15:0]data_in_R_47_I,
    input [15:0]data_in_R_47_Q,
    input [15:0]data_in_R_48_I,
    input [15:0]data_in_R_48_Q,
    input [15:0]data_in_R_49_I,
    input [15:0]data_in_R_49_Q,
    input [15:0]data_in_R_50_I,
    input [15:0]data_in_R_50_Q,
    input [15:0]data_in_R_51_I,
    input [15:0]data_in_R_51_Q,
    input [15:0]data_in_R_52_I,
    input [15:0]data_in_R_52_Q,
    input [15:0]data_in_R_53_I,
    input [15:0]data_in_R_53_Q,
    input [15:0]data_in_R_54_I,
    input [15:0]data_in_R_54_Q,
    input [15:0]data_in_R_55_I,
    input [15:0]data_in_R_55_Q,
    input [15:0]data_in_R_56_I,
    input [15:0]data_in_R_56_Q,
    input [15:0]data_in_R_57_I,
    input [15:0]data_in_R_57_Q,
    input [15:0]data_in_R_58_I,
    input [15:0]data_in_R_58_Q,
    input [15:0]data_in_R_59_I,
    input [15:0]data_in_R_59_Q,
    input [15:0]data_in_R_60_I,
    input [15:0]data_in_R_60_Q,
    input [15:0]data_in_R_61_I,
    input [15:0]data_in_R_61_Q,
    input [15:0]data_in_R_62_I,
    input [15:0]data_in_R_62_Q,
    input [15:0]data_in_R_63_I,
    input [15:0]data_in_R_63_Q,
    input [15:0]data_in_R_64_I,
    input [15:0]data_in_R_64_Q,
    input [15:0]data_in_R_65_I,
    input [15:0]data_in_R_65_Q,
    input [15:0]data_in_R_66_I,
    input [15:0]data_in_R_66_Q,
    input [15:0]data_in_R_67_I,
    input [15:0]data_in_R_67_Q,
    input [15:0]data_in_R_68_I,
    input [15:0]data_in_R_68_Q,
    input [15:0]data_in_R_69_I,
    input [15:0]data_in_R_69_Q,
    input [15:0]data_in_R_70_I,
    input [15:0]data_in_R_70_Q,
    

    
    output [15:0]add_L_1_35_I,
    output [15:0]add_L_1_35_Q,
    output [15:0]add_R_1_35_I,
    output [15:0]add_R_1_35_Q,
    output [15:0]add_L_36_70_I,
    output [15:0]add_L_36_70_Q,
    output [15:0]add_R_36_70_I,
    output [15:0]add_R_36_70_Q,
    output dataout_valid
    );
    wire dataout_valid_1;
    wire [15:0]add_L_1_35_I_2 ;
    wire [15:0]add_L_1_35_Q_2 ;
    wire [15:0]add_R_1_35_I_2 ;
    wire [15:0]add_R_1_35_Q_2 ;
    wire [15:0]add_L_36_70_I_2;
    wire [15:0]add_L_36_70_Q_2;
    wire [15:0]add_R_36_70_I_2;
    wire [15:0]add_R_36_70_Q_2; 
    
    wire [21:0]add_L_1_35_I_1 ;
    wire [21:0]add_L_1_35_Q_1 ;
    wire [21:0]add_R_1_35_I_1 ;
    wire [21:0]add_R_1_35_Q_1 ;
    wire [21:0]add_L_36_70_I_1;
    wire [21:0]add_L_36_70_Q_1;
    wire [21:0]add_R_36_70_I_1;
    wire [21:0]add_R_36_70_Q_1; 
add_1_35  add_l_1_35( 
  .clk(clk),     
     .data_in_I1 (data_in_L_1_I ),
     .data_in_Q1 (data_in_L_1_Q ),
     .data_in_I2 (data_in_L_2_I ),
     .data_in_Q2 (data_in_L_2_Q ),
     .data_in_I3 (data_in_L_3_I ),
     .data_in_Q3 (data_in_L_3_Q ),
     .data_in_I4 (data_in_L_4_I ),
     .data_in_Q4 (data_in_L_4_Q ),
     .data_in_I5 (data_in_L_5_I ),
     .data_in_Q5 (data_in_L_5_Q ),
     .data_in_I6 (data_in_L_6_I ),
     .data_in_Q6 (data_in_L_6_Q ),
     .data_in_I7 (data_in_L_7_I ),
     .data_in_Q7 (data_in_L_7_Q ),
     .data_in_I8 (data_in_L_8_I ),
     .data_in_Q8 (data_in_L_8_Q ),
     .data_in_I9 (data_in_L_9_I ),
     .data_in_Q9 (data_in_L_9_Q ),
     .data_in_I10(data_in_L_10_I),
     .data_in_Q10(data_in_L_10_Q),
     .data_in_I11(data_in_L_11_I),
     .data_in_Q11(data_in_L_11_Q),
     .data_in_I12(data_in_L_12_I),
     .data_in_Q12(data_in_L_12_Q),
     .data_in_I13(data_in_L_13_I),
     .data_in_Q13(data_in_L_13_Q),
     .data_in_I14(data_in_L_14_I),
     .data_in_Q14(data_in_L_14_Q),
     .data_in_I15(data_in_L_15_I),
     .data_in_Q15(data_in_L_15_Q),
     .data_in_I16(data_in_L_16_I),
     .data_in_Q16(data_in_L_16_Q),
     .data_in_I17(data_in_L_17_I),
     .data_in_Q17(data_in_L_17_Q),
     .data_in_I18(data_in_L_18_I),
     .data_in_Q18(data_in_L_18_Q),
     .data_in_I19(data_in_L_19_I),
     .data_in_Q19(data_in_L_19_Q),
     .data_in_I20(data_in_L_20_I),
     .data_in_Q20(data_in_L_20_Q),
     .data_in_I21(data_in_L_21_I),
     .data_in_Q21(data_in_L_21_Q),
     .data_in_I22(data_in_L_22_I),
     .data_in_Q22(data_in_L_22_Q),
     .data_in_I23(data_in_L_23_I),
     .data_in_Q23(data_in_L_23_Q),
     .data_in_I24(data_in_L_24_I),
     .data_in_Q24(data_in_L_24_Q),
     .data_in_I25(data_in_L_25_I),
     .data_in_Q25(data_in_L_25_Q),
     .data_in_I26(data_in_L_26_I),
     .data_in_Q26(data_in_L_26_Q),
     .data_in_I27(data_in_L_27_I),
     .data_in_Q27(data_in_L_27_Q),
     .data_in_I28(data_in_L_28_I),
     .data_in_Q28(data_in_L_28_Q),
     .data_in_I29(data_in_L_29_I),
     .data_in_Q29(data_in_L_29_Q),
     .data_in_I30(data_in_L_30_I),
     .data_in_Q30(data_in_L_30_Q),
     .data_in_I31(data_in_L_31_I),
     .data_in_Q31(data_in_L_31_Q),
     .data_in_I32(data_in_L_32_I),
     .data_in_Q32(data_in_L_32_Q),
     .data_in_I33(data_in_L_33_I),
     .data_in_Q33(data_in_L_33_Q),
     .data_in_I34(data_in_L_34_I),
     .data_in_Q34(data_in_L_34_Q),
     .data_in_I35(data_in_L_35_I),
     .data_in_Q35(data_in_L_35_Q),
     .data_in_valid(data_in_valid),
     .sum_1_35_I(add_L_1_35_I_1),
     .sum_1_35_Q(add_L_1_35_Q_1),
     .data_out_valid(dataout_valid_1)  
       
) ;   

add_1_35  add_r_1_35(    
  .clk(clk),  
     .data_in_I1 (data_in_R_1_I ),
     .data_in_Q1 (data_in_R_1_Q ),
     .data_in_I2 (data_in_R_2_I ),
     .data_in_Q2 (data_in_R_2_Q ),
     .data_in_I3 (data_in_R_3_I ),
     .data_in_Q3 (data_in_R_3_Q ),
     .data_in_I4 (data_in_R_4_I ),
     .data_in_Q4 (data_in_R_4_Q ),
     .data_in_I5 (data_in_R_5_I ),
     .data_in_Q5 (data_in_R_5_Q ),
     .data_in_I6 (data_in_R_6_I ),
     .data_in_Q6 (data_in_R_6_Q ),
     .data_in_I7 (data_in_R_7_I ),
     .data_in_Q7 (data_in_R_7_Q ),
     .data_in_I8 (data_in_R_8_I ),
     .data_in_Q8 (data_in_R_8_Q ),
     .data_in_I9 (data_in_R_9_I ),
     .data_in_Q9 (data_in_R_9_Q ),
     .data_in_I10(data_in_R_10_I),
     .data_in_Q10(data_in_R_10_Q),
     .data_in_I11(data_in_R_11_I),
     .data_in_Q11(data_in_R_11_Q),
     .data_in_I12(data_in_R_12_I),
     .data_in_Q12(data_in_R_12_Q),
     .data_in_I13(data_in_R_13_I),
     .data_in_Q13(data_in_R_13_Q),
     .data_in_I14(data_in_R_14_I),
     .data_in_Q14(data_in_R_14_Q),
     .data_in_I15(data_in_R_15_I),
     .data_in_Q15(data_in_R_15_Q),
     .data_in_I16(data_in_R_16_I),
     .data_in_Q16(data_in_R_16_Q),
     .data_in_I17(data_in_R_17_I),
     .data_in_Q17(data_in_R_17_Q),
     .data_in_I18(data_in_R_18_I),
     .data_in_Q18(data_in_R_18_Q),
     .data_in_I19(data_in_R_19_I),
     .data_in_Q19(data_in_R_19_Q),
     .data_in_I20(data_in_R_20_I),
     .data_in_Q20(data_in_R_20_Q),
     .data_in_I21(data_in_R_21_I),
     .data_in_Q21(data_in_R_21_Q),
     .data_in_I22(data_in_R_22_I),
     .data_in_Q22(data_in_R_22_Q),
     .data_in_I23(data_in_R_23_I),
     .data_in_Q23(data_in_R_23_Q),
     .data_in_I24(data_in_R_24_I),
     .data_in_Q24(data_in_R_24_Q),
     .data_in_I25(data_in_R_25_I),
     .data_in_Q25(data_in_R_25_Q),
     .data_in_I26(data_in_R_26_I),
     .data_in_Q26(data_in_R_26_Q),
     .data_in_I27(data_in_R_27_I),
     .data_in_Q27(data_in_R_27_Q),
     .data_in_I28(data_in_R_28_I),
     .data_in_Q28(data_in_R_28_Q),
     .data_in_I29(data_in_R_29_I),
     .data_in_Q29(data_in_R_29_Q),
     .data_in_I30(data_in_R_30_I),
     .data_in_Q30(data_in_R_30_Q),
     .data_in_I31(data_in_R_31_I),
     .data_in_Q31(data_in_R_31_Q),
     .data_in_I32(data_in_R_32_I),
     .data_in_Q32(data_in_R_32_Q),
     .data_in_I33(data_in_R_33_I),
     .data_in_Q33(data_in_R_33_Q),
     .data_in_I34(data_in_R_34_I),
     .data_in_Q34(data_in_R_34_Q),
     .data_in_I35(data_in_R_35_I),
     .data_in_Q35(data_in_R_35_Q),
     .data_in_valid(data_in_valid),
     .sum_1_35_I(add_R_1_35_I_1),
     .sum_1_35_Q(add_R_1_35_Q_1),
     .data_out_valid()  
       
) ;  
add_1_35  add_l_36_70(  
  .clk(clk),    
     .data_in_I1 (data_in_L_36_I),
     .data_in_Q1 (data_in_L_36_Q),
     .data_in_I2 (data_in_L_37_I),
     .data_in_Q2 (data_in_L_37_Q),
     .data_in_I3 (data_in_L_38_I),
     .data_in_Q3 (data_in_L_38_Q),
     .data_in_I4 (data_in_L_39_I),
     .data_in_Q4 (data_in_L_39_Q),
     .data_in_I5 (data_in_L_40_I),
     .data_in_Q5 (data_in_L_40_Q),
     .data_in_I6 (data_in_L_41_I),
     .data_in_Q6 (data_in_L_41_Q),
     .data_in_I7 (data_in_L_42_I),
     .data_in_Q7 (data_in_L_42_Q),
     .data_in_I8 (data_in_L_43_I),
     .data_in_Q8 (data_in_L_43_Q),
     .data_in_I9 (data_in_L_44_I),
     .data_in_Q9 (data_in_L_44_Q),
     .data_in_I10(data_in_L_45_I),
     .data_in_Q10(data_in_L_45_Q),
     .data_in_I11(data_in_L_46_I),
     .data_in_Q11(data_in_L_46_Q),
     .data_in_I12(data_in_L_47_I),
     .data_in_Q12(data_in_L_47_Q),
     .data_in_I13(data_in_L_48_I),
     .data_in_Q13(data_in_L_48_Q),
     .data_in_I14(data_in_L_49_I),
     .data_in_Q14(data_in_L_49_Q),
     .data_in_I15(data_in_L_50_I),
     .data_in_Q15(data_in_L_50_Q),
     .data_in_I16(data_in_L_51_I),
     .data_in_Q16(data_in_L_51_Q),
     .data_in_I17(data_in_L_52_I),
     .data_in_Q17(data_in_L_52_Q),
     .data_in_I18(data_in_L_53_I),
     .data_in_Q18(data_in_L_53_Q),
     .data_in_I19(data_in_L_54_I),
     .data_in_Q19(data_in_L_54_Q),
     .data_in_I20(data_in_L_55_I),
     .data_in_Q20(data_in_L_55_Q),
     .data_in_I21(data_in_L_56_I),
     .data_in_Q21(data_in_L_56_Q),
     .data_in_I22(data_in_L_57_I),
     .data_in_Q22(data_in_L_57_Q),
     .data_in_I23(data_in_L_58_I),
     .data_in_Q23(data_in_L_58_Q),
     .data_in_I24(data_in_L_59_I),
     .data_in_Q24(data_in_L_59_Q),
     .data_in_I25(data_in_L_60_I),
     .data_in_Q25(data_in_L_60_Q),
     .data_in_I26(data_in_L_61_I),
     .data_in_Q26(data_in_L_61_Q),
     .data_in_I27(data_in_L_62_I),
     .data_in_Q27(data_in_L_62_Q),
     .data_in_I28(data_in_L_63_I),
     .data_in_Q28(data_in_L_63_Q),
     .data_in_I29(data_in_L_64_I),
     .data_in_Q29(data_in_L_64_Q),
     .data_in_I30(data_in_L_65_I),
     .data_in_Q30(data_in_L_65_Q),
     .data_in_I31(data_in_L_66_I),
     .data_in_Q31(data_in_L_66_Q),
     .data_in_I32(data_in_L_67_I),
     .data_in_Q32(data_in_L_67_Q),
     .data_in_I33(data_in_L_68_I),
     .data_in_Q33(data_in_L_68_Q),
     .data_in_I34(data_in_L_69_I),
     .data_in_Q34(data_in_L_69_Q),
     .data_in_I35(data_in_L_70_I),
     .data_in_Q35(data_in_L_70_Q),
     .data_in_valid(data_in_valid),
     .sum_1_35_I(add_L_36_70_I_1),
     .sum_1_35_Q(add_L_36_70_Q_1),
     .data_out_valid()  
       
) ;  

add_1_35  add_r_36_70(    
  .clk(clk),  
     .data_in_I1 (data_in_R_36_I),
     .data_in_Q1 (data_in_R_36_Q),
     .data_in_I2 (data_in_R_37_I),
     .data_in_Q2 (data_in_R_37_Q),
     .data_in_I3 (data_in_R_38_I),
     .data_in_Q3 (data_in_R_38_Q),
     .data_in_I4 (data_in_R_39_I),
     .data_in_Q4 (data_in_R_39_Q),
     .data_in_I5 (data_in_R_40_I),
     .data_in_Q5 (data_in_R_40_Q),
     .data_in_I6 (data_in_R_41_I),
     .data_in_Q6 (data_in_R_41_Q),
     .data_in_I7 (data_in_R_42_I),
     .data_in_Q7 (data_in_R_42_Q),
     .data_in_I8 (data_in_R_43_I),
     .data_in_Q8 (data_in_R_43_Q),
     .data_in_I9 (data_in_R_44_I),
     .data_in_Q9 (data_in_R_44_Q),
     .data_in_I10(data_in_R_45_I),
     .data_in_Q10(data_in_R_45_Q),
     .data_in_I11(data_in_R_46_I),
     .data_in_Q11(data_in_R_46_Q),
     .data_in_I12(data_in_R_47_I),
     .data_in_Q12(data_in_R_47_Q),
     .data_in_I13(data_in_R_48_I),
     .data_in_Q13(data_in_R_48_Q),
     .data_in_I14(data_in_R_49_I),
     .data_in_Q14(data_in_R_49_Q),
     .data_in_I15(data_in_R_50_I),
     .data_in_Q15(data_in_R_50_Q),
     .data_in_I16(data_in_R_51_I),
     .data_in_Q16(data_in_R_51_Q),
     .data_in_I17(data_in_R_52_I),
     .data_in_Q17(data_in_R_52_Q),
     .data_in_I18(data_in_R_53_I),
     .data_in_Q18(data_in_R_53_Q),
     .data_in_I19(data_in_R_54_I),
     .data_in_Q19(data_in_R_54_Q),
     .data_in_I20(data_in_R_55_I),
     .data_in_Q20(data_in_R_55_Q),
     .data_in_I21(data_in_R_56_I),
     .data_in_Q21(data_in_R_56_Q),
     .data_in_I22(data_in_R_57_I),
     .data_in_Q22(data_in_R_57_Q),
     .data_in_I23(data_in_R_58_I),
     .data_in_Q23(data_in_R_58_Q),
     .data_in_I24(data_in_R_59_I),
     .data_in_Q24(data_in_R_59_Q),
     .data_in_I25(data_in_R_60_I),
     .data_in_Q25(data_in_R_60_Q),
     .data_in_I26(data_in_R_61_I),
     .data_in_Q26(data_in_R_61_Q),
     .data_in_I27(data_in_R_62_I),
     .data_in_Q27(data_in_R_62_Q),
     .data_in_I28(data_in_R_63_I),
     .data_in_Q28(data_in_R_63_Q),
     .data_in_I29(data_in_R_64_I),
     .data_in_Q29(data_in_R_64_Q),
     .data_in_I30(data_in_R_65_I),
     .data_in_Q30(data_in_R_65_Q),
     .data_in_I31(data_in_R_66_I),
     .data_in_Q31(data_in_R_66_Q),
     .data_in_I32(data_in_R_67_I),
     .data_in_Q32(data_in_R_67_Q),
     .data_in_I33(data_in_R_68_I),
     .data_in_Q33(data_in_R_68_Q),
     .data_in_I34(data_in_R_69_I),
     .data_in_Q34(data_in_R_69_Q),
     .data_in_I35(data_in_R_70_I),
     .data_in_Q35(data_in_R_70_Q),
     .data_in_valid(data_in_valid),
     .sum_1_35_I(add_R_36_70_I_1),
     .sum_1_35_Q(add_R_36_70_Q_1),
     .data_out_valid()  
       
) ;  
wire dataout_valid_2;
wire [2:0]cut_ctl;
vio_add_cut vio_add_cut_1 (
  .clk(clk),                // input wire clk
  .probe_out0(cut_ctl)  // output wire [2 : 0] probe_out0
);
cut_add  #(.LEN(22))
                 add_cut_1(
    .clk(clk),
    .data_i(add_L_1_35_I_1),
    .data_q(add_L_1_35_Q_1),
    .in_valid(dataout_valid_1),
    .cut_ctl(cut_ctl),
    
    .data_out_i(add_L_1_35_I_2),
    .data_out_q(add_L_1_35_Q_2),
    .out_valid(dataout_valid_2)
    );
    
cut_add  #(.LEN(22))
                 add_cut_2(
    .clk(clk),
    .data_i(add_R_1_35_I_1),
    .data_q(add_R_1_35_Q_1),
    .in_valid(dataout_valid_1),
    .cut_ctl(cut_ctl),
    
    .data_out_i(add_R_1_35_I_2),
    .data_out_q(add_R_1_35_Q_2),
    .out_valid()
    );
    
cut_add  #(.LEN(22))
                add_cut_3(
    .clk(clk),
    .data_i(add_L_36_70_I_1),
    .data_q(add_L_36_70_Q_1),
    .in_valid(dataout_valid_1),
    .cut_ctl(cut_ctl),
    
    .data_out_i(add_L_36_70_I_2),
    .data_out_q(add_L_36_70_Q_2),
    .out_valid()
    );
    
cut_add  #(.LEN(22))
                 add_cut_4(
    .clk(clk),
    .data_i(add_R_36_70_I_1),
    .data_q(add_R_36_70_Q_1),
    .in_valid(dataout_valid_1),
    .cut_ctl(cut_ctl),
    
    .data_out_i(add_R_36_70_I_2),
    .data_out_q(add_R_36_70_Q_2),
    .out_valid()
    );
assign dataout_valid = dataout_valid_2;
assign add_L_1_35_I  = add_L_1_35_I_2 ;
assign add_L_1_35_Q  = add_L_1_35_Q_2 ;
assign add_R_1_35_I  = add_R_1_35_I_2 ;
assign add_R_1_35_Q  = add_R_1_35_Q_2 ;
assign add_L_36_70_I = add_L_36_70_I_2;
assign add_L_36_70_Q = add_L_36_70_Q_2;
assign add_R_36_70_I = add_R_36_70_I_2;
assign add_R_36_70_Q = add_R_36_70_Q_2;

ila_aaaa ila_aaa (
	.clk(clk), // input wire clk


	.probe0(data_in_valid), // input wire [0:0]  probe0  
	.probe1(dataout_valid_1), // input wire [0:0]  probe1 
	.probe2(dataout_valid_2), // input wire [0:0]  probe2 
	.probe3(dataout_valid), // input wire [0:0]  probe3 
	.probe4(data_in_L_1_I), // input wire [15:0]  probe4 
	.probe5(data_in_L_1_Q), // input wire [15:0]  probe5 
	.probe6(add_L_1_35_I_1), // input wire [21:0]  probe6 
	.probe7(add_L_1_35_Q_1), // input wire [21:0]  probe7 
	.probe8(add_L_1_35_I), // input wire [15:0]  probe8 
	.probe9(add_L_1_35_Q), // input wire [15:0]  probe9
    .probe10(add_R_1_35_I), // input wire [15:0]  probe10 
	.probe11(add_R_1_35_Q), // input wire [15:0]  probe11 
	.probe12(add_L_36_70_Q), // input wire [15:0]  probe12 
	.probe13(add_L_36_70_Q), // input wire [15:0]  probe13 
	.probe14(add_R_36_70_Q), // input wire [15:0]  probe14 
	.probe15(add_R_36_70_Q) // input wire [15:0]  probe15
	
	
	
	
);
endmodule
