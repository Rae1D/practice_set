`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/09/10 11:33:35
// Design Name: 
// Module Name: dbf_fangwei
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module dbf_fangwei(
    input clk_120m,
    input [15:0] dataI,
    input [15:0] dataQ,
    input data_in_valid,                        ////////////******************
    
    input [3:0]fpga_gpio,
    
    output [15:0]add_out_1_24_I,
    output [15:0]add_out_1_24_Q,
    output [15:0]add_out_25_48_I,
    output [15:0]add_out_25_48_Q,
    output data_out_valid   

    );
    wire [2:0]fw_cut_ctl ;
    wire [15:0] A;
    reg phase_data_valid = 1;          /////////////************
   vio_fangwei_cut vio_fangwei_cut_1 (
  .clk(clk_120m),                // input wire clk
  .probe_out0(fw_cut_ctl)  // output wire [2 : 0] probe_out0
); 
    wire [15:0] A_fw;
    reg  fangwei_rst = 1;

//    vio_FW tt (
//      .clk(clk_120m),                // input wire clk
//      .probe_in0(fpga_gpio[0]),    // input wire [0 : 0] probe_in0
//      .probe_out0(fangwei_rst),  // output wire [0 : 0] probe_out0
//      .probe_out1(A_fw),  // output wire [0 : 0] probe_out0
//      .probe_out2(fw_cut_ctl)  // output wire [0 : 0] probe_out0
//    );
//    assign A = A_fw;
///////////////////////////////////////
    reg [15:0]A_1  = 16'b0010111101100010;
    reg [15:0]A_2  = 16'b0011000000100000; 
    reg [15:0]A_3  = 16'b0011000110011001;
    reg [15:0]A_4  = 16'b0011001111001000;
    reg [15:0]A_5  = 16'b0011011010100100;
    reg [15:0]A_6  = 16'b0011101000100011;
    reg [15:0]A_7  = 16'b0011111000110100;
    reg [15:0]A_8  = 16'b0100001011000101;
    reg [15:0]A_9  = 16'b0100011110111110;
    reg [15:0]A_10 = 16'b0100110100000101;
    reg [15:0]A_11 = 16'b0101001001111101;
    reg [15:0]A_12 = 16'b0101100000001000;
    reg [15:0]A_13 = 16'b0101110110000110;
    reg [15:0]A_14 = 16'b0110001011011011;
    reg [15:0]A_15 = 16'b0110011111101011;
    reg [15:0]A_16 = 16'b0110110010011111;
    reg [15:0]A_17 = 16'b0111000011100100;
    reg [15:0]A_18 = 16'b0111010010101011;
    reg [15:0]A_19 = 16'b0111011111101100;
    reg [15:0]A_20 = 16'b0111101010100010;
    reg [15:0]A_21 = 16'b0111110011001010;
    reg [15:0]A_22 = 16'b0111111001100110;
    reg [15:0]A_23 = 16'b0111111101110111;
    reg [15:0]A_24 = 16'b0111111111111111;
    reg [15:0]A_25 = 16'b0111111111111111;
    reg [15:0]A_26 = 16'b0111111101110111;
    reg [15:0]A_27 = 16'b0111111001100110;
    reg [15:0]A_28 = 16'b0111110011001010;
    reg [15:0]A_29 = 16'b0111101010100010;
    reg [15:0]A_30 = 16'b0111011111101100;
    reg [15:0]A_31 = 16'b0111010010101011;
    reg [15:0]A_32 = 16'b0111000011100100;
    reg [15:0]A_33 = 16'b0110110010011111;
    reg [15:0]A_34 = 16'b0110011111101011;
    reg [15:0]A_35 = 16'b0110001011011011;
    reg [15:0]A_36 = 16'b0101110110000110;
    reg [15:0]A_37 = 16'b0101100000001000;
    reg [15:0]A_38 = 16'b0101001001111101;
    reg [15:0]A_39 = 16'b0100110100000101;
    reg [15:0]A_40 = 16'b0100011110111110;
    reg [15:0]A_41 = 16'b0100001011000101;
    reg [15:0]A_42 = 16'b0011111000110100;
    reg [15:0]A_43 = 16'b0011101000100011;
    reg [15:0]A_44 = 16'b0011011010100100;
    reg [15:0]A_45 = 16'b0011001111001000;
    reg [15:0]A_46 = 16'b0011000110011001;
    reg [15:0]A_47 = 16'b0011000000100000;
    reg [15:0]A_48 = 16'b0010111101100010;
   

reg   [15:0]ph_real_1   ;
reg   [15:0]ph_real_2   ;
reg   [15:0]ph_real_3   ;
reg   [15:0]ph_real_4   ;
reg   [15:0]ph_real_5   ;
reg   [15:0]ph_real_6   ;
reg   [15:0]ph_real_7   ;
reg   [15:0]ph_real_8   ;
reg   [15:0]ph_real_9   ;
reg   [15:0]ph_real_10   ;
reg   [15:0]ph_real_11   ;
reg   [15:0]ph_real_12   ;
reg   [15:0]ph_real_13   ;
reg   [15:0]ph_real_14   ;
reg   [15:0]ph_real_15  ;
reg   [15:0]ph_real_16   ;
reg   [15:0]ph_real_17   ;
reg   [15:0]ph_real_18   ;
reg   [15:0]ph_real_19   ;
reg   [15:0]ph_real_20   ;
reg   [15:0]ph_real_21   ;   
reg   [15:0]ph_real_22   ;
reg   [15:0]ph_real_23   ;
reg   [15:0]ph_real_24   ;
reg   [15:0]ph_real_25   ;
reg   [15:0]ph_real_26   ;
reg   [15:0]ph_real_27   ;
reg   [15:0]ph_real_28   ;   
reg   [15:0]ph_real_29    ;
reg   [15:0]ph_real_30   ;
reg   [15:0]ph_real_31   ;
reg   [15:0]ph_real_32   ;
reg   [15:0]ph_real_33   ;
reg   [15:0]ph_real_34   ;
reg   [15:0]ph_real_35   ;
reg   [15:0]ph_real_36   ;
reg   [15:0]ph_real_37   ;
reg   [15:0]ph_real_38   ;
reg   [15:0]ph_real_39   ;
reg   [15:0]ph_real_40   ;
reg   [15:0]ph_real_41   ;
reg   [15:0]ph_real_42   ;
reg   [15:0]ph_real_43  ;
reg   [15:0]ph_real_44   ;
reg   [15:0]ph_real_45   ;
reg   [15:0]ph_real_46   ;
reg   [15:0]ph_real_47   ;
reg   [15:0]ph_real_48   ;

                 
reg   [15:0]ph_image_1  ;
reg   [15:0]ph_image_2  ;
reg   [15:0]ph_image_3  ;
reg   [15:0]ph_image_4  ;
reg   [15:0]ph_image_5  ;
reg   [15:0]ph_image_6  ;
reg   [15:0]ph_image_7  ;
reg   [15:0]ph_image_8  ;
reg   [15:0]ph_image_9  ;
reg   [15:0]ph_image_10 ;
reg   [15:0]ph_image_11 ;
reg   [15:0]ph_image_12 ;
reg   [15:0]ph_image_13 ;
reg   [15:0]ph_image_14 ;
reg   [15:0]ph_image_15 ;
reg   [15:0]ph_image_16 ;
reg   [15:0]ph_image_17 ;
reg   [15:0]ph_image_18 ;
reg   [15:0]ph_image_19 ;
reg   [15:0]ph_image_20 ;
reg   [15:0]ph_image_21 ;
reg   [15:0]ph_image_22 ;
reg   [15:0]ph_image_23 ;
reg   [15:0]ph_image_24 ;
reg   [15:0]ph_image_25 ;
reg   [15:0]ph_image_26 ;
reg   [15:0]ph_image_27 ;
reg   [15:0]ph_image_28 ;
reg   [15:0]ph_image_29 ;
reg   [15:0]ph_image_30 ;
reg   [15:0]ph_image_31 ;
reg   [15:0]ph_image_32 ;
reg   [15:0]ph_image_33 ;
reg   [15:0]ph_image_34 ;
reg   [15:0]ph_image_35 ;
reg   [15:0]ph_image_36 ;
reg   [15:0]ph_image_37 ;
reg   [15:0]ph_image_38 ;
reg   [15:0]ph_image_39 ;
reg   [15:0]ph_image_40 ;
reg   [15:0]ph_image_41 ;
reg   [15:0]ph_image_42 ;
reg   [15:0]ph_image_43 ;
reg   [15:0]ph_image_44 ;
reg   [15:0]ph_image_45 ;
reg   [15:0]ph_image_46 ;
reg   [15:0]ph_image_47 ;
reg   [15:0]ph_image_48 ;
/////////////////////////////////////////////////////////////////  
wire [4:0]fw_fcode;
vio_fw_fcode fw_f (
  .clk(clk_120m),                // input wire clk
  .probe_out0(fw_fcode)  // output wire [4 : 0] probe_out0
);

always@(posedge clk_120m)
begin
    case(fw_fcode)
    0: begin
        if(fpga_gpio == 4'b0000)   ///////频点0----目标波达方向0.25°----接收方位波束指向0°  
       begin
       ph_real_1  <=  16'b0011111111111111;
       ph_real_2  <=  16'b0011111111111101;
       ph_real_3  <=  16'b0011111111110110;
       ph_real_4  <=  16'b0011111111101100;
       ph_real_5  <=  16'b0011111111011101;
       ph_real_6  <=  16'b0011111111001010;
       ph_real_7  <=  16'b0011111110110010;
       ph_real_8  <=  16'b0011111110010110;
       ph_real_9  <=  16'b0011111101110110;
       ph_real_10  <= 16'b0011111101010010;
       ph_real_11  <= 16'b0011111100101010;
       ph_real_12  <= 16'b0011111011111101;
       ph_real_13  <= 16'b0011111011001100;
       ph_real_14  <= 16'b0011111010010111;
       ph_real_15  <= 16'b0011111001011110;
       ph_real_16  <= 16'b0011111000100000;
       ph_real_17  <= 16'b0011110111011111;
       ph_real_18  <= 16'b0011110110011001;
       ph_real_19  <= 16'b0011110101001111;
       ph_real_20  <= 16'b0011110100000001;
       ph_real_21  <= 16'b0011110010101111;
       ph_real_22  <= 16'b0011110001011001;
       ph_real_23  <= 16'b0011101111111111;
       ph_real_24  <= 16'b0011101110100001;
       ph_real_25  <= 16'b0011101100111111;
       ph_real_26  <= 16'b0011101011011001;
       ph_real_27  <= 16'b0011101001101111;
       ph_real_28  <= 16'b0011101000000001;
       ph_real_29  <= 16'b0011100110001111;
       ph_real_30  <= 16'b0011100100011001;
       ph_real_31  <= 16'b0011100010100000;
       ph_real_32  <= 16'b0011100000100011;
       ph_real_33  <= 16'b0011011110100010;
       ph_real_34  <= 16'b0011011100011101;
       ph_real_35  <= 16'b0011011010010101;
       ph_real_36  <= 16'b0011011000001001;
       ph_real_37  <= 16'b0011010101111001;
       ph_real_38  <= 16'b0011010011100110;
       ph_real_39  <= 16'b0011010001001111;
       ph_real_40  <= 16'b0011001110110101;
       ph_real_41  <= 16'b0011001100010111;
       ph_real_42  <= 16'b0011001001110110;
       ph_real_43  <= 16'b0011000111010001;
       ph_real_44  <= 16'b0011000100101010;
       ph_real_45  <= 16'b0011000001111110;
       ph_real_46  <= 16'b0010111111010000;
       ph_real_47  <= 16'b0010111100011111;
       ph_real_48  <= 16'b0010111001101010;
       
      ph_image_1 =  16'b0000000000000000;
      ph_image_2 =  16'b0000000100001000;
      ph_image_3 =  16'b0000001000010001; 
      ph_image_4 =  16'b0000001100011001;
      ph_image_5 =  16'b0000010000100010;
      ph_image_6 =  16'b0000010100101010;
      ph_image_7 =  16'b0000011000110001;
      ph_image_8 =  16'b0000011100111000;
      ph_image_9 =  16'b0000100000111111;
      ph_image_10<= 16'b0000100101000101;
      ph_image_11<= 16'b0000101001001011;
      ph_image_12<= 16'b0000101101010000;
      ph_image_13<= 16'b0000110001010100;
      ph_image_14<= 16'b0000110101010111;
      ph_image_15<= 16'b0000111001011010;
      ph_image_16<= 16'b0000111101011011;
      ph_image_17<= 16'b0001000001011100;
      ph_image_18<= 16'b0001000101011011;
      ph_image_19<= 16'b0001001001011001;
      ph_image_20<= 16'b0001001101010110;
      ph_image_21<= 16'b0001010001010010;
      ph_image_22<= 16'b0001010101001100;
      ph_image_23<= 16'b0001011001000101;
      ph_image_24<= 16'b0001011100111101;
      ph_image_25<= 16'b0001100000110010;
      ph_image_26<= 16'b0001100100100111;
      ph_image_27<= 16'b0001101000011001;
      ph_image_28<= 16'b0001101100001010;
      ph_image_29<= 16'b0001101111111001;
      ph_image_30<= 16'b0001110011100110;
      ph_image_31<= 16'b0001110111010001;
      ph_image_32<= 16'b0001111010111011;
      ph_image_33<= 16'b0001111110100010;
      ph_image_34<= 16'b0010000010000111;
      ph_image_35<= 16'b0010000101101010; 
      ph_image_36<= 16'b0010001001001010;
      ph_image_37<= 16'b0010001100101001;
      ph_image_38<= 16'b0010010000000101;
      ph_image_39<= 16'b0010010011011110;
      ph_image_40<= 16'b0010010110110101;
      ph_image_41<= 16'b0010011010001010;
      ph_image_42<= 16'b0010011101011100;
      ph_image_43<= 16'b0010100000101011;
      ph_image_44<= 16'b0010100011111000;
      ph_image_45<= 16'b0010100111000010;
      ph_image_46<= 16'b0010101010001001;
      ph_image_47<= 16'b0010101101001110;
      ph_image_48<= 16'b0010110000001111;
      
       end
       else if(fpga_gpio == 4'b0001)    ///////频点0----目标波达方向-0.25°----接收方位波束指向0°  
       begin
       ph_real_1  <=  16'b0011111111111111;
       ph_real_2  <=  16'b0011111111111101;
       ph_real_3  <=  16'b0011111111110110; 
       ph_real_4  <=  16'b0011111111101100;
       ph_real_5  <=  16'b0011111111011101;
       ph_real_6  <=  16'b0011111111001010;
       ph_real_7  <=  16'b0011111110110010;
       ph_real_8  <=  16'b0011111110010110;
       ph_real_9  <=  16'b0011111101110110;
       ph_real_10  <= 16'b0011111101010010;
       ph_real_11  <= 16'b0011111100101010;
       ph_real_12  <= 16'b0011111011111101;
       ph_real_13  <= 16'b0011111011001100;
       ph_real_14  <= 16'b0011111010010111;
       ph_real_15  <= 16'b0011111001011110;
       ph_real_16  <= 16'b0011111000100000;
       ph_real_17  <= 16'b0011110111011111;
       ph_real_18  <= 16'b0011110110011001;
       ph_real_19  <= 16'b0011110101001111;
       ph_real_20  <= 16'b0011110100000001;
       ph_real_21  <= 16'b0011110010101111;
       ph_real_22  <= 16'b0011110001011001;
       ph_real_23  <= 16'b0011101111111111;
       ph_real_24  <= 16'b0011101110100001;
       ph_real_25  <= 16'b0011101100111111;
       ph_real_26  <= 16'b0011101011011001;
       ph_real_27  <= 16'b0011101001101111;
       ph_real_28  <= 16'b0011101000000001;
       ph_real_29  <= 16'b0011100110001111;
       ph_real_30  <= 16'b0011100100011001;
       ph_real_31  <= 16'b0011100010100000;
       ph_real_32  <= 16'b0011100000100011;
       ph_real_33  <= 16'b0011011110100010;
       ph_real_34  <= 16'b0011011100011101;
       ph_real_35  <= 16'b0011011010010101; 
       ph_real_36  <= 16'b0011011000001001;
       ph_real_37  <= 16'b0011010101111001;
       ph_real_38  <= 16'b0011010011100110;
       ph_real_39  <= 16'b0011010001001111;
       ph_real_40  <= 16'b0011001110110101;
       ph_real_41  <= 16'b0011001100010111;
       ph_real_42  <= 16'b0011001001110110;
       ph_real_43  <= 16'b0011000111010001;
       ph_real_44  <= 16'b0011000100101010;
       ph_real_45  <= 16'b0011000001111110;
       ph_real_46  <= 16'b0010111111010000;
       ph_real_47  <= 16'b0010111100011111;
       ph_real_48  <= 16'b0010111001101010;
       
      ph_image_1 =  16'b0000000000000000;
      ph_image_2 =  16'b1111111011110111;
      ph_image_3 =  16'b1111110111101111; 
      ph_image_4 =  16'b1111110011100110;
      ph_image_5 =  16'b1111101111011110;
      ph_image_6 =  16'b1111101011010110;
      ph_image_7 =  16'b1111100111001110;
      ph_image_8 =  16'b1111100011000111;
      ph_image_9 =  16'b1111011111000000;
      ph_image_10<= 16'b1111011010111010;
      ph_image_11<= 16'b1111010110110100;
      ph_image_12<= 16'b1111010010110000;
      ph_image_13<= 16'b1111001110101011;
      ph_image_14<= 16'b1111001010101000;
      ph_image_15<= 16'b1111000110100110;
      ph_image_16<= 16'b1111000010100100;
      ph_image_17<= 16'b1110111110100100;
      ph_image_18<= 16'b1110111010100100;
      ph_image_19<= 16'b1110110110100110;
      ph_image_20<= 16'b1110110010101001;
      ph_image_21<= 16'b1110101110101110;
      ph_image_22<= 16'b1110101010110011;
      ph_image_23<= 16'b1110100110111010;
      ph_image_24<= 16'b1110100011000011;
      ph_image_25<= 16'b1110011111001101;
      ph_image_26<= 16'b1110011011011001;
      ph_image_27<= 16'b1110010111100110;
      ph_image_28<= 16'b1110010011110101;
      ph_image_29<= 16'b1110010000000110;
      ph_image_30<= 16'b1110001100011001;
      ph_image_31<= 16'b1110001000101110;
      ph_image_32<= 16'b1110000101000101;
      ph_image_33<= 16'b1110000001011110;
      ph_image_34<= 16'b1101111101111001;
      ph_image_35<= 16'b1101111010010110; 
      ph_image_36<= 16'b1101110110110101;
      ph_image_37<= 16'b1101110011010111;
      ph_image_38<= 16'b1101101111111011;
      ph_image_39<= 16'b1101101100100001;
      ph_image_40<= 16'b1101101001001010;
      ph_image_41<= 16'b1101100101110110;
      ph_image_42<= 16'b1101100010100100;
      ph_image_43<= 16'b1101011111010100;
      ph_image_44<= 16'b1101011100000111;
      ph_image_45<= 16'b1101011000111101;
      ph_image_46<= 16'b1101010101110110;
      ph_image_47<= 16'b1101010010110010;
      ph_image_48<= 16'b1101001111110001;
       end
       
       
    ////////////////////////////////////////////
       else if(fpga_gpio == 4'b0010)   ///////频点0----目标波达方向0.75°----接收方位波束指向0°  
       begin 
       ph_real_1  <=  16'b0011111111111111;
       ph_real_2  <=  16'b0011111111101100;
       ph_real_3  <=  16'b0011111110110010; 
       ph_real_4  <=  16'b0011111101010010;
       ph_real_5  <=  16'b0011111011001100;
       ph_real_6  <=  16'b0011111000100000;
       ph_real_7  <=  16'b0011110101001111;
       ph_real_8  <=  16'b0011110001011001;
       ph_real_9  <=  16'b0011101100111111;
       ph_real_10  <= 16'b0011101000000001;
       ph_real_11  <= 16'b0011100010100000;
       ph_real_12  <= 16'b0011011100011101;
       ph_real_13  <= 16'b0011010101111001;
       ph_real_14  <= 16'b0011001110110101;
       ph_real_15  <= 16'b0011000111010010;
       ph_real_16  <= 16'b0010111111010000;
       ph_real_17  <= 16'b0010110110110010;
       ph_real_18  <= 16'b0010101101111001;
       ph_real_19  <= 16'b0010100100100101;
       ph_real_20  <= 16'b0010011010111001;
       ph_real_21  <= 16'b0010010000110101;
       ph_real_22  <= 16'b0010000110011100;
       ph_real_23  <= 16'b0001111011101110;
       ph_real_24  <= 16'b0001110000101110;
       ph_real_25  <= 16'b0001100101011101;
       ph_real_26  <= 16'b0001011001111101;
       ph_real_27  <= 16'b0001001110001111;
       ph_real_28  <= 16'b0001000010010101;
       ph_real_29  <= 16'b0000110110010001;
       ph_real_30  <= 16'b0000101010000110;
       ph_real_31  <= 16'b0000011101110011;
       ph_real_32  <= 16'b0000010001011101;
       ph_real_33  <= 16'b0000000101000100;
       ph_real_34  <= 16'b1111111000101010;
       ph_real_35  <= 16'b1111101100010001; 
       ph_real_36  <= 16'b1111011111111011;
       ph_real_37  <= 16'b1111010011101010;
       ph_real_38  <= 16'b1111000111100000;
       ph_real_39  <= 16'b1110111011011110;
       ph_real_40  <= 16'b1110101111100110;
       ph_real_41  <= 16'b1110100011111010;
       ph_real_42  <= 16'b1110011000011101;
       ph_real_43  <= 16'b1110001101001110;
       ph_real_44  <= 16'b1110000010010010;
       ph_real_45  <= 16'b1101110111101000;
       ph_real_46  <= 16'b1101101101010010;
       ph_real_47  <= 16'b1101100011010011;
       ph_real_48  <= 16'b1101011001101011;
       
      ph_image_1 =  16'b0000000000000000;
      ph_image_2 =  16'b0000001100011001;
      ph_image_3 =  16'b0000011000110001; 
      ph_image_4 =  16'b0000100101000101;
      ph_image_5 =  16'b0000110001010100;
      ph_image_6 =  16'b0000111101011011;
      ph_image_7 =  16'b0001001001011001;
      ph_image_8 =  16'b0001010101001100;
      ph_image_9 =  16'b0001100000110010;
      ph_image_10<= 16'b0001101100001010;
      ph_image_11<= 16'b0001110111010001;
      ph_image_12<= 16'b0010000010000111;
      ph_image_13<= 16'b0010001100101000;
      ph_image_14<= 16'b0010010110110101;
      ph_image_15<= 16'b0010100000101011;
      ph_image_16<= 16'b0010101010001001;
      ph_image_17<= 16'b0010110011001101;
      ph_image_18<= 16'b0010111011110111;
      ph_image_19<= 16'b0011000100000100;
      ph_image_20<= 16'b0011001011110011;
      ph_image_21<= 16'b0011010011000100;
      ph_image_22<= 16'b0011011001110110;
      ph_image_23<= 16'b0011100000000110;
      ph_image_24<= 16'b0011100101110101;
      ph_image_25<= 16'b0011101011000001;
      ph_image_26<= 16'b0011101111101010;
      ph_image_27<= 16'b0011110011101111;
      ph_image_28<= 16'b0011110111001111;
      ph_image_29<= 16'b0011111010001010;
      ph_image_30<= 16'b0011111100100000;
      ph_image_31<= 16'b0011111110010000;
      ph_image_32<= 16'b0011111111011001;
      ph_image_33<= 16'b0011111111111100;
      ph_image_34<= 16'b0011111111111000;
      ph_image_35<= 16'b0011111111001110; 
      ph_image_36<= 16'b0011111101111110;
      ph_image_37<= 16'b0011111100000111;
      ph_image_38<= 16'b0011111001101011;
      ph_image_39<= 16'b0011110110101001;
      ph_image_40<= 16'b0011110011000010;
      ph_image_41<= 16'b0011101110110110;
      ph_image_42<= 16'b0011101010000111;
      ph_image_43<= 16'b0011100100110100;
      ph_image_44<= 16'b0011011110111111;
      ph_image_45<= 16'b0011011000101000;
      ph_image_46<= 16'b0011010001110001;
      ph_image_47<= 16'b0011001010011010;
      ph_image_48<= 16'b0011000010100101;
       end
       else if(fpga_gpio == 4'b0011)   ///////频点0----目标波达方向-0.75°----接收方位波束指向0°  
       begin
       ph_real_1  <=  16'b0011111111111111;
       ph_real_2  <=  16'b0011111111101100;
       ph_real_3  <=  16'b0011111110110010; 
       ph_real_4  <=  16'b0011111101010010;
       ph_real_5  <=  16'b0011111011001100;
       ph_real_6  <=  16'b0011111000100000;
       ph_real_7  <=  16'b0011110101001111;
       ph_real_8  <=  16'b0011110001011001;
       ph_real_9  <=  16'b0011101100111111;
       ph_real_10  <= 16'b0011101000000001;
       ph_real_11  <= 16'b0011100010100000;
       ph_real_12  <= 16'b0011011100011101;
       ph_real_13  <= 16'b0011010101111001;
       ph_real_14  <= 16'b0011001110110101;
       ph_real_15  <= 16'b0011000111010010;
       ph_real_16  <= 16'b0010111111010000;
       ph_real_17  <= 16'b0010110110110010;
       ph_real_18  <= 16'b0010101101111001;
       ph_real_19  <= 16'b0010100100100101;
       ph_real_20  <= 16'b0010011010111001;
       ph_real_21  <= 16'b0010010000110101;
       ph_real_22  <= 16'b0010000110011100;
       ph_real_23  <= 16'b0001111011101110;
       ph_real_24  <= 16'b0001110000101110;
       ph_real_25  <= 16'b0001100101011101;
       ph_real_26  <= 16'b0001011001111101;
       ph_real_27  <= 16'b0001001110001111;
       ph_real_28  <= 16'b0001000010010101;
       ph_real_29  <= 16'b0000110110010001;
       ph_real_30  <= 16'b0000101010000110;
       ph_real_31  <= 16'b0000011101110011;
       ph_real_32  <= 16'b0000010001011101;
       ph_real_33  <= 16'b0000000101000100;
       ph_real_34  <= 16'b1111111000101010;
       ph_real_35  <= 16'b1111101100010001; 
       ph_real_36  <= 16'b1111011111111011;
       ph_real_37  <= 16'b1111010011101010;
       ph_real_38  <= 16'b1111000111100000;
       ph_real_39  <= 16'b1110111011011110;
       ph_real_40  <= 16'b1110101111100110;
       ph_real_41  <= 16'b1110100011111010;
       ph_real_42  <= 16'b1110011000011101;
       ph_real_43  <= 16'b1110001101001110;
       ph_real_44  <= 16'b1110000010010010;
       ph_real_45  <= 16'b1101110111101000;
       ph_real_46  <= 16'b1101101101010010;
       ph_real_47  <= 16'b1101100011010011;
       ph_real_48  <= 16'b1101011001101011;
       
      ph_image_1 =  16'b0000000000000000;
      ph_image_2 =  16'b1111110011100110;
      ph_image_3 =  16'b1111100111001110; 
      ph_image_4 =  16'b1111011010111010;
      ph_image_5 =  16'b1111001110101011;
      ph_image_6 =  16'b1111000010100100;
      ph_image_7 =  16'b1110110110100110;
      ph_image_8 =  16'b1110101010110011;
      ph_image_9 =  16'b1110011111001101;
      ph_image_10<= 16'b1110010011110110;
      ph_image_11<= 16'b1110001000101110;
      ph_image_12<= 16'b1101111101111001;
      ph_image_13<= 16'b1101110011010111;
      ph_image_14<= 16'b1101101001001010;
      ph_image_15<= 16'b1101011111010100;
      ph_image_16<= 16'b1101010101110111;
      ph_image_17<= 16'b1101001100110010;
      ph_image_18<= 16'b1101000100001001;
      ph_image_19<= 16'b1100111011111100;
      ph_image_20<= 16'b1100110100001100;
      ph_image_21<= 16'b1100101100111011;
      ph_image_22<= 16'b1100100110001010;
      ph_image_23<= 16'b1100011111111001;
      ph_image_24<= 16'b1100011010001011;
      ph_image_25<= 16'b1100010100111110;
      ph_image_26<= 16'b1100010000010101;
      ph_image_27<= 16'b1100001100010000;
      ph_image_28<= 16'b1100001000110000;
      ph_image_29<= 16'b1100000101110101;
      ph_image_30<= 16'b1100000011100000;
      ph_image_31<= 16'b1100000001110000;
      ph_image_32<= 16'b1100000000100111;
      ph_image_33<= 16'b1100000000000100;
      ph_image_34<= 16'b1100000000000111;
      ph_image_35<= 16'b1100000000110001; 
      ph_image_36<= 16'b1100000010000010;
      ph_image_37<= 16'b1100000011111000;
      ph_image_38<= 16'b1100000110010101;
      ph_image_39<= 16'b1100001001010111;
      ph_image_40<= 16'b1100001100111110;
      ph_image_41<= 16'b1100010001001001;
      ph_image_42<= 16'b1100010101111001;
      ph_image_43<= 16'b1100011011001011;
      ph_image_44<= 16'b1100100001000001;
      ph_image_45<= 16'b1100100111010111;
      ph_image_46<= 16'b1100101110001110;
      ph_image_47<= 16'b1100110101100101;
      ph_image_48<= 16'b1100111101011010;
       end
    ////////////////////////////////////////////
       else if(fpga_gpio == 4'b0100)   ///////频点0----目标波达方向1.5°----接收方位波束指向0°  
       begin 
       ph_real_1  <=  16'b0011111111111111;
       ph_real_2  <=  16'b0011111110110010;
       ph_real_3  <=  16'b0011111011001100; 
       ph_real_4  <=  16'b0011110101001111;
       ph_real_5  <=  16'b0011101100111111;
       ph_real_6  <=  16'b0011100010100000;
       ph_real_7  <=  16'b0011010101111001;
       ph_real_8  <=  16'b0011000111010010;
       ph_real_9  <=  16'b0010110110110011;
       ph_real_10  <= 16'b0010100100100110;
       ph_real_11  <= 16'b0010010000110110;
       ph_real_12  <= 16'b0001111011110000;
       ph_real_13  <= 16'b0001100101011111;
       ph_real_14  <= 16'b0001001110010000;
       ph_real_15  <= 16'b0000110110010011;
       ph_real_16  <= 16'b0000011101110101;
       ph_real_17  <= 16'b0000000101000110;
       ph_real_18  <= 16'b1111101100010011;
       ph_real_19  <= 16'b1111010011101100;
       ph_real_20  <= 16'b1110111011100000;
       ph_real_21  <= 16'b1110100011111101;
       ph_real_22  <= 16'b1110001101010001;
       ph_real_23  <= 16'b1101110111101010;
       ph_real_24  <= 16'b1101100011010101;
       ph_real_25  <= 16'b1101010000011110;
       ph_real_26  <= 16'b1100111111010001;
       ph_real_27  <= 16'b1100101111110111;
       ph_real_28  <= 16'b1100100010011011;
       ph_real_29  <= 16'b1100010111000011;
       ph_real_30  <= 16'b1100001101111000;
       ph_real_31  <= 16'b1100000110111110;
       ph_real_32  <= 16'b1100000010011001;
       ph_real_33  <= 16'b1100000000001101;
       ph_real_34  <= 16'b1100000000011011;
       ph_real_35  <= 16'b1100000011000010; 
       ph_real_36  <= 16'b1100001000000010;
       ph_real_37  <= 16'b1100001111010110;
       ph_real_38  <= 16'b1100011000111011;
       ph_real_39  <= 16'b1100100100101011;
       ph_real_40  <= 16'b1100110010011110;
       ph_real_41  <= 16'b1101000010001101;
       ph_real_42  <= 16'b1101010011101110;
       ph_real_43  <= 16'b1101100110110111;
       ph_real_44  <= 16'b1101111011011011;
       ph_real_45  <= 16'b1110010001001111;
       ph_real_46  <= 16'b1110101000000110;
       ph_real_47  <= 16'b1110111111110010;
       ph_real_48  <= 16'b1111011000000100;
      
      ph_image_1 =  16'b0000000000000000;
      ph_image_2 =  16'b0000011000110001;
      ph_image_3 =  16'b0000110001010100; 
      ph_image_4 =  16'b0001001001011001;
      ph_image_5 =  16'b0001100000110010;
      ph_image_6 =  16'b0001110111010001;
      ph_image_7 =  16'b0010001100101000;
      ph_image_8 =  16'b0010100000101010;
      ph_image_9 =  16'b0010110011001100;
      ph_image_10<= 16'b0011000100000011;
      ph_image_11<= 16'b0011010011000100;
      ph_image_12<= 16'b0011100000000101;
      ph_image_13<= 16'b0011101011000001;
      ph_image_14<= 16'b0011110011101111;
      ph_image_15<= 16'b0011111010001010;
      ph_image_16<= 16'b0011111110001111;
      ph_image_17<= 16'b0011111111111100;
      ph_image_18<= 16'b0011111111001110;
      ph_image_19<= 16'b0011111100001000;
      ph_image_20<= 16'b0011110110101010;
      ph_image_21<= 16'b0011101110110111;
      ph_image_22<= 16'b0011100100110101;
      ph_image_23<= 16'b0011011000101010;
      ph_image_24<= 16'b0011001010011100;
      ph_image_25<= 16'b0010111010010101;
      ph_image_26<= 16'b0010101000011110;
      ph_image_27<= 16'b0010010101000010;
      ph_image_28<= 16'b0010000000001100;
      ph_image_29<= 16'b0001101010001001;
      ph_image_30<= 16'b0001010011000110;
      ph_image_31<= 16'b0000111011010001;
      ph_image_32<= 16'b0000100010111001;
      ph_image_33<= 16'b0000001010001100;
      ph_image_34<= 16'b1111110001011001;
      ph_image_35<= 16'b1111011000101110; 
      ph_image_36<= 16'b1111000000011011;
      ph_image_37<= 16'b1110101000101110;
      ph_image_38<= 16'b1110010001110110;
      ph_image_39<= 16'b1101111100000000;
      ph_image_40<= 16'b1101100111011001;
      ph_image_41<= 16'b1101010100001110;
      ph_image_42<= 16'b1101000010101010;
      ph_image_43<= 16'b1100110010111000;
      ph_image_44<= 16'b1100100101000001;
      ph_image_45<= 16'b1100011001001101;
      ph_image_46<= 16'b1100001111100101;
      ph_image_47<= 16'b1100001000001100;
      ph_image_48<= 16'b1100000011001001;
       end
       else if(fpga_gpio == 4'b0101)   ///////频点0----目标波达方向-1.5°----接收方位波束指向0°  
       begin
       ph_real_1  <=  16'b0011111111111111;
       ph_real_2  <=  16'b0011111110110010;
       ph_real_3  <=  16'b0011111011001100; 
       ph_real_4  <=  16'b0011110101001111;
       ph_real_5  <=  16'b0011101100111111;
       ph_real_6  <=  16'b0011100010100000;
       ph_real_7  <=  16'b0011010101111001;
       ph_real_8  <=  16'b0011000111010010;
       ph_real_9  <=  16'b0010110110110011;
       ph_real_10  <= 16'b0010100100100110;
       ph_real_11  <= 16'b0010010000110110;
       ph_real_12  <= 16'b0001111011110000;
       ph_real_13  <= 16'b0001100101011111;
       ph_real_14  <= 16'b0001001110010000;
       ph_real_15  <= 16'b0000110110010011;
       ph_real_16  <= 16'b0000011101110101;
       ph_real_17  <= 16'b0000000101000110;
       ph_real_18  <= 16'b1111101100010011;
       ph_real_19  <= 16'b1111010011101100;
       ph_real_20  <= 16'b1110111011100000;
       ph_real_21  <= 16'b1110100011111101;
       ph_real_22  <= 16'b1110001101010001;
       ph_real_23  <= 16'b1101110111101010;
       ph_real_24  <= 16'b1101100011010101;
       ph_real_25  <= 16'b1101010000011110;
       ph_real_26  <= 16'b1100111111010001;
       ph_real_27  <= 16'b1100101111110111;
       ph_real_28  <= 16'b1100100010011011;
       ph_real_29  <= 16'b1100010111000011;
       ph_real_30  <= 16'b1100001101111000;
       ph_real_31  <= 16'b1100000110111110;
       ph_real_32  <= 16'b1100000010011001;
       ph_real_33  <= 16'b1100000000001101;
       ph_real_34  <= 16'b1100000000011011;
       ph_real_35  <= 16'b1100000011000010; 
       ph_real_36  <= 16'b1100001000000010;
       ph_real_37  <= 16'b1100001111010110;
       ph_real_38  <= 16'b1100011000111011;
       ph_real_39  <= 16'b1100100100101011;
       ph_real_40  <= 16'b1100110010011110;
       ph_real_41  <= 16'b1101000010001101;
       ph_real_42  <= 16'b1101010011101110;
       ph_real_43  <= 16'b1101100110110111;
       ph_real_44  <= 16'b1101111011011011;
       ph_real_45  <= 16'b1110010001001111;
       ph_real_46  <= 16'b1110101000000110;
       ph_real_47  <= 16'b1110111111110010;
       ph_real_48  <= 16'b1111011000000100;
       
      ph_image_1 =  16'b0000000000000000;
      ph_image_2 =  16'b1111100111001110;
      ph_image_3 =  16'b1111001110101100; 
      ph_image_4 =  16'b1110110110100111;
      ph_image_5 =  16'b1110011111001110;
      ph_image_6 =  16'b1110001000101111;
      ph_image_7 =  16'b1101110011011000;
      ph_image_8 =  16'b1101011111010101;
      ph_image_9 =  16'b1101001100110011;
      ph_image_10<= 16'b1100111011111101;
      ph_image_11<= 16'b1100101100111100;
      ph_image_12<= 16'b1100011111111010;
      ph_image_13<= 16'b1100010100111111;
      ph_image_14<= 16'b1100001100010001;
      ph_image_15<= 16'b1100000101110101;
      ph_image_16<= 16'b1100000001110000;
      ph_image_17<= 16'b1100000000000100;
      ph_image_18<= 16'b1100000000110001;
      ph_image_19<= 16'b1100000011111000;
      ph_image_20<= 16'b1100001001010110;
      ph_image_21<= 16'b1100010001001000;
      ph_image_22<= 16'b1100011011001010;
      ph_image_23<= 16'b1100100111010110;
      ph_image_24<= 16'b1100110101100011;
      ph_image_25<= 16'b1101000101101010;
      ph_image_26<= 16'b1101010111100010;
      ph_image_27<= 16'b1101101010111110;
      ph_image_28<= 16'b1101111111110100;
      ph_image_29<= 16'b1110010101110111;
      ph_image_30<= 16'b1110101100111010;
      ph_image_31<= 16'b1111000100101110;
      ph_image_32<= 16'b1111011101000111;
      ph_image_33<= 16'b1111110101110100;
      ph_image_34<= 16'b0000001110100111;
      ph_image_35<= 16'b0000100111010001; 
      ph_image_36<= 16'b0000111111100100;
      ph_image_37<= 16'b0001010111010001;
      ph_image_38<= 16'b0001101110001001;
      ph_image_39<= 16'b0010000100000000;
      ph_image_40<= 16'b0010011000100110;
      ph_image_41<= 16'b0010101011110010;
      ph_image_42<= 16'b0010111101010110;
      ph_image_43<= 16'b0011001101001000;
      ph_image_44<= 16'b0011011010111111;
      ph_image_45<= 16'b0011100110110010;
      ph_image_46<= 16'b0011110000011011;
      ph_image_47<= 16'b0011110111110011;
      ph_image_48<= 16'b0011111100110110;
       end
    ////////////////////////////////////////////
       else if(fpga_gpio == 4'b0110)   ///////频点0----目标波达方向3.5°----接收方位波束指向0°  
       begin 
       ph_real_1  <=  16'b0011111111111111;
       ph_real_2  <=  16'b0011111001011110;
       ph_real_3  <=  16'b0011100110010001; 
       ph_real_4  <=  16'b0011000111010110;
       ph_real_5  <=  16'b0010011110010001;
       ph_real_6  <=  16'b0001101101001010;
       ph_real_7  <=  16'b0000110110011110;
       ph_real_8  <=  16'b1111111101000010;
       ph_real_9  <=  16'b1111000011101111;
       ph_real_10  <= 16'b1110001101100000;
       ph_real_11  <= 16'b1101011101000110;
       ph_real_12  <= 16'b1100110100111111;
       ph_real_13  <= 16'b1100010111001101;
       ph_real_14  <= 16'b1100000101010000;
       ph_real_15  <= 16'b1100000000000101;
       ph_real_16  <= 16'b1100000111111011;
       ph_real_17  <= 16'b1100011100011001;
       ph_real_18  <= 16'b1100111100011100;
       ph_real_19  <= 16'b1101100110011011;
       ph_real_20  <= 16'b1110011000010000;
       ph_real_21  <= 16'b1111001111010101;
       ph_real_22  <= 16'b0000001000111001;
       ph_real_23  <= 16'b0001000010000001;
       ph_real_24  <= 16'b0001110111110001;
       ph_real_25  <= 16'b0010100111011100;
       ph_real_26  <= 16'b0011001110100101;
       ph_real_27  <= 16'b0011101011001101;
       ph_real_28  <= 16'b0011111011110111;
       ph_real_29  <= 16'b0011111111101101;
       ph_real_30  <= 16'b0011110110100011;
       ph_real_31  <= 16'b0011100000110101;
       ph_real_32  <= 16'b0010111111101011;
       ph_real_33  <= 16'b0010010100110001;
       ph_real_34  <= 16'b0001100010010011;
       ph_real_35  <= 16'b0000101010110100; 
       ph_real_36  <= 16'b1111110001001011;
       ph_real_37  <= 16'b1110111000010001;
       ph_real_38  <= 16'b1110000011000001;
       ph_real_39  <= 16'b1101010100000111;
       ph_real_40  <= 16'b1100101101111110;
       ph_real_41  <= 16'b1100010010100001;
       ph_real_42  <= 16'b1100000011001001;
       ph_real_43  <= 16'b1100000000101000;
       ph_real_44  <= 16'b1100001011000111;
       ph_real_45  <= 16'b1100100010000100;
       ph_real_46  <= 16'b1101000100010011;
       ph_real_47  <= 16'b1101110000000110;
       ph_real_48  <= 16'b1110100011001101;
       
      ph_image_1 =  16'b0000000000000000;
      ph_image_2 =  16'b0000111001011000;
      ph_image_3 =  16'b0001101111110101; 
      ph_image_4 =  16'b0010100000100110;
      ph_image_5 =  16'b0011001001001100;
      ph_image_6 =  16'b0011100111100011;
      ph_image_7 =  16'b0011111010001000;
      ph_image_8 =  16'b0011111111111110;
      ph_image_9 =  16'b0011111000110011;
      ph_image_10<= 16'b0011100100111101;
      ph_image_11<= 16'b0011000101011110;
      ph_image_12<= 16'b0010011011111011;
      ph_image_13<= 16'b0001101010011101;
      ph_image_14<= 16'b0000110011100100;
      ph_image_15<= 16'b1111111010000100;
      ph_image_16<= 16'b1111000000110111;
      ph_image_17<= 16'b1110001010110111;
      ph_image_18<= 16'b1101011010110100;
      ph_image_19<= 16'b1100110011001100;
      ph_image_20<= 16'b1100010101111111;
      ph_image_21<= 16'b1100000100101011;
      ph_image_22<= 16'b1100000000001010;
      ph_image_23<= 16'b1100001000101011;
      ph_image_24<= 16'b1100011101110000;
      ph_image_25<= 16'b1100111110010111;
      ph_image_26<= 16'b1101101000110100;
      ph_image_27<= 16'b1110011010111110;
      ph_image_28<= 16'b1111010010010000;
      ph_image_29<= 16'b0000001011110111;
      ph_image_30<= 16'b0001000100111000;
      ph_image_31<= 16'b0001111010011001;
      ph_image_32<= 16'b0010101001101010;
      ph_image_33<= 16'b0011010000010100;
      ph_image_34<= 16'b0011101100010111;
      ph_image_35<= 16'b0011111100011000; 
      ph_image_36<= 16'b0011111111100011;
      ph_image_37<= 16'b0011110101101111;
      ph_image_38<= 16'b0011011111011001;
      ph_image_39<= 16'b0010111101101101;
      ph_image_40<= 16'b0010010010010110;
      ph_image_41<= 16'b0001011111100011;
      ph_image_42<= 16'b0000100111111001;
      ph_image_43<= 16'b1111101110001101;
      ph_image_44<= 16'b1110110101011011;
      ph_image_45<= 16'b1110000000011011;
      ph_image_46<= 16'b1101010001111011;
      ph_image_47<= 16'b1100101100010010;
      ph_image_48<= 16'b1100010001011011;
       end
       
       else if(fpga_gpio == 4'b0111)   ///////频点0----目标波达方向-3.5°----接收方位波束指向0°  
       begin
       ph_real_1  <=  16'b0011111111111111;
       ph_real_2  <=  16'b0011111001011110;
       ph_real_3  <=  16'b0011100110010001; 
       ph_real_4  <=  16'b0011000111010110;
       ph_real_5  <=  16'b0010011110010001;
       ph_real_6  <=  16'b0001101101001010;
       ph_real_7  <=  16'b0000110110011110;
       ph_real_8  <=  16'b1111111101000010;
       ph_real_9  <=  16'b1111000011101111;
       ph_real_10  <= 16'b1110001101100000;
       ph_real_11  <= 16'b1101011101000110;
       ph_real_12  <= 16'b1100110100111111;
       ph_real_13  <= 16'b1100010111001101;
       ph_real_14  <= 16'b1100000101010000;
       ph_real_15  <= 16'b1100000000000101;
       ph_real_16  <= 16'b1100000111111011;
       ph_real_17  <= 16'b1100011100011001;
       ph_real_18  <= 16'b1100111100011100;
       ph_real_19  <= 16'b1101100110011011;
       ph_real_20  <= 16'b1110011000010000;
       ph_real_21  <= 16'b1111001111010101;
       ph_real_22  <= 16'b0000001000111001;
       ph_real_23  <= 16'b0001000010000001;
       ph_real_24  <= 16'b0001110111110001;
       ph_real_25  <= 16'b0010100111011100;
       ph_real_26  <= 16'b0011001110100101;
       ph_real_27  <= 16'b0011101011001101;
       ph_real_28  <= 16'b0011111011110111;
       ph_real_29  <= 16'b0011111111101101;
       ph_real_30  <= 16'b0011110110100011;
       ph_real_31  <= 16'b0011100000110101;
       ph_real_32  <= 16'b0010111111101011;
       ph_real_33  <= 16'b0010010100110001;
       ph_real_34  <= 16'b0001100010010011;
       ph_real_35  <= 16'b0000101010110100; 
       ph_real_36  <= 16'b1111110001001011;
       ph_real_37  <= 16'b1110111000010001;
       ph_real_38  <= 16'b1110000011000001;
       ph_real_39  <= 16'b1101010100000111;
       ph_real_40  <= 16'b1100101101111110;
       ph_real_41  <= 16'b1100010010100001;
       ph_real_42  <= 16'b1100000011001001;
       ph_real_43  <= 16'b1100000000101000;
       ph_real_44  <= 16'b1100001011000111;
       ph_real_45  <= 16'b1100100010000100;
       ph_real_46  <= 16'b1101000100010011;
       ph_real_47  <= 16'b1101110000000110;
       ph_real_48  <= 16'b1110100011001101;
       
      ph_image_1 =  16'b0000000000000000;
      ph_image_2 =  16'b1111000110101000;
      ph_image_3 =  16'b1110010000001011; 
      ph_image_4 =  16'b1101011111011010;
      ph_image_5 =  16'b1100110110110011;
      ph_image_6 =  16'b1100011000011101;
      ph_image_7 =  16'b1100000101111000;
      ph_image_8 =  16'b1100000000000010;
      ph_image_9 =  16'b1100000111001101;
      ph_image_10<= 16'b1100011011000011;
      ph_image_11<= 16'b1100111010100010;
      ph_image_12<= 16'b1101100100000100;
      ph_image_13<= 16'b1110010101100010;
      ph_image_14<= 16'b1111001100011011;
      ph_image_15<= 16'b0000000101111011;
      ph_image_16<= 16'b0000111111001001;
      ph_image_17<= 16'b0001110101001001;
      ph_image_18<= 16'b0010100101001011;
      ph_image_19<= 16'b0011001100110011;
      ph_image_20<= 16'b0011101010000001;
      ph_image_21<= 16'b0011111011010100;
      ph_image_22<= 16'b0011111111110101;
      ph_image_23<= 16'b0011110111010101;
      ph_image_24<= 16'b0011100010001111;
      ph_image_25<= 16'b0011000001101000;
      ph_image_26<= 16'b0010010111001011;
      ph_image_27<= 16'b0001100101000010;
      ph_image_28<= 16'b0000101101101111;
      ph_image_29<= 16'b1111110100001000;
      ph_image_30<= 16'b1110111011000111;
      ph_image_31<= 16'b1110000101100111;
      ph_image_32<= 16'b1101010110010101;
      ph_image_33<= 16'b1100101111101100;
      ph_image_34<= 16'b1100010011101001;
      ph_image_35<= 16'b1100000011100111; 
      ph_image_36<= 16'b1100000000011100;
      ph_image_37<= 16'b1100001010010001;
      ph_image_38<= 16'b1100100000100110;
      ph_image_39<= 16'b1101000010010011;
      ph_image_40<= 16'b1101101101101001;
      ph_image_41<= 16'b1110100000011100;
      ph_image_42<= 16'b1111011000000111;
      ph_image_43<= 16'b0000010001110010;
      ph_image_44<= 16'b0001001010100101;
      ph_image_45<= 16'b0001111111100100;
      ph_image_46<= 16'b0010101110000100;
      ph_image_47<= 16'b0011010011101101;
      ph_image_48<= 16'b0011101110100101;
       end
   
      
    ////////////////////////////////////////////
       else 
       begin
       ph_real_1  <=  16'b0011111111111111;
       ph_real_2  <=  16'b0011111111111111;
       ph_real_3  <=  16'b0011111111111111; 
       ph_real_4  <=  16'b0011111111111111;
       ph_real_5  <=  16'b0011111111111111;
       ph_real_6  <=  16'b0011111111111111;
       ph_real_7  <=  16'b0011111111111111;
       ph_real_8  <=  16'b0011111111111111;
       ph_real_9  <=  16'b0011111111111111;
       ph_real_10  <= 16'b0011111111111111;
       ph_real_11  <= 16'b0011111111111111;
       ph_real_12  <= 16'b0011111111111111;
       ph_real_13  <= 16'b0011111111111111;
       ph_real_14  <= 16'b0011111111111111;
       ph_real_15  <= 16'b0011111111111111;
       ph_real_16  <= 16'b0011111111111111;
       ph_real_17  <= 16'b0011111111111111;
       ph_real_18  <= 16'b0011111111111111;
       ph_real_19  <= 16'b0011111111111111;
       ph_real_20  <= 16'b0011111111111111;
       ph_real_21  <= 16'b0011111111111111;
       ph_real_22  <= 16'b0011111111111111;
       ph_real_23  <= 16'b0011111111111111;
       ph_real_24  <= 16'b0011111111111111;
       ph_real_25  <= 16'b0011111111111111;
       ph_real_26  <= 16'b0011111111111111;
       ph_real_27  <= 16'b0011111111111111;
       ph_real_28  <= 16'b0011111111111111;
       ph_real_29  <= 16'b0011111111111111;
       ph_real_30  <= 16'b0011111111111111;
       ph_real_31  <= 16'b0011111111111111;
       ph_real_32  <= 16'b0011111111111111;
       ph_real_33  <= 16'b0011111111111111;
       ph_real_34  <= 16'b0011111111111111;
       ph_real_35  <= 16'b0011111111111111; 
       ph_real_36  <= 16'b0011111111111111;
       ph_real_37  <= 16'b0011111111111111;
       ph_real_38  <= 16'b0011111111111111;
       ph_real_39  <= 16'b0011111111111111;
       ph_real_40  <= 16'b0011111111111111;
       ph_real_41  <= 16'b0011111111111111;
       ph_real_42  <= 16'b0011111111111111;
       ph_real_43  <= 16'b0011111111111111;
       ph_real_44  <= 16'b0011111111111111;
       ph_real_45  <= 16'b0011111111111111;
       ph_real_46  <= 16'b0011111111111111;
       ph_real_47  <= 16'b0011111111111111;
       ph_real_48  <= 16'b0011111111111111;
       
      ph_image_1 =  16'b0000000000000000;
      ph_image_2 =  16'b0000000000000000;
      ph_image_3 =  16'b0000000000000000; 
      ph_image_4 =  16'b0000000000000000;
      ph_image_5 =  16'b0000000000000000;
      ph_image_6 =  16'b0000000000000000;
      ph_image_7 =  16'b0000000000000000;
      ph_image_8 =  16'b0000000000000000;
      ph_image_9 =  16'b0000000000000000;
      ph_image_10<= 16'b0000000000000000;
      ph_image_11<= 16'b0000000000000000;
      ph_image_12<= 16'b0000000000000000;
      ph_image_13<= 16'b0000000000000000;
      ph_image_14<= 16'b0000000000000000;
      ph_image_15<= 16'b0000000000000000;
      ph_image_16<= 16'b0000000000000000;
      ph_image_17<= 16'b0000000000000000;
      ph_image_18<= 16'b0000000000000000;
      ph_image_19<= 16'b0000000000000000;
      ph_image_20<= 16'b0000000000000000;
      ph_image_21<= 16'b0000000000000000;
      ph_image_22<= 16'b0000000000000000;
      ph_image_23<= 16'b0000000000000000;
      ph_image_24<= 16'b0000000000000000;
      ph_image_25<= 16'b0000000000000000;
      ph_image_26<= 16'b0000000000000000;
      ph_image_27<= 16'b0000000000000000;
      ph_image_28<= 16'b0000000000000000;
      ph_image_29<= 16'b0000000000000000;
      ph_image_30<= 16'b0000000000000000;
      ph_image_31<= 16'b0000000000000000;
      ph_image_32<= 16'b0000000000000000;
      ph_image_33<= 16'b0000000000000000;
      ph_image_34<= 16'b0000000000000000;
      ph_image_35<= 16'b0000000000000000; 
      ph_image_36<= 16'b0000000000000000;
      ph_image_37<= 16'b0000000000000000;
      ph_image_38<= 16'b0000000000000000;
      ph_image_39<= 16'b0000000000000000;
      ph_image_40<= 16'b0000000000000000;
      ph_image_41<= 16'b0000000000000000;
      ph_image_42<= 16'b0000000000000000;
      ph_image_43<= 16'b0000000000000000;
      ph_image_44<= 16'b0000000000000000;
      ph_image_45<= 16'b0000000000000000;
      ph_image_46<= 16'b0000000000000000;
      ph_image_47<= 16'b0000000000000000;
      ph_image_48<= 16'b0000000000000000;
       end
    ////////////////////////////////////////////
        end
   
     
    default:          
       begin
       ph_real_1  <=  16'b0000000000000000;
       ph_real_2  <=  16'b0000000000000000;
       ph_real_3  <=  16'b0000000000000000; 
       ph_real_4  <=  16'b0000000000000000;
       ph_real_5  <=  16'b0000000000000000;
       ph_real_6  <=  16'b0000000000000000;
       ph_real_7  <=  16'b0000000000000000;
       ph_real_8  <=  16'b0000000000000000;
       ph_real_9  <=  16'b0000000000000000;
       ph_real_10  <= 16'b0000000000000000;
       ph_real_11  <= 16'b0000000000000000;
       ph_real_12  <= 16'b0000000000000000;
       ph_real_13  <= 16'b0000000000000000;
       ph_real_14  <= 16'b0000000000000000;
       ph_real_15  <= 16'b0000000000000000;
       ph_real_16  <= 16'b0000000000000000;
       ph_real_17  <= 16'b0000000000000000;
       ph_real_18  <= 16'b0000000000000000;
       ph_real_19  <= 16'b0000000000000000;
       ph_real_20  <= 16'b0000000000000000;
       ph_real_21  <= 16'b0000000000000000;
       ph_real_22  <= 16'b0000000000000000;
       ph_real_23  <= 16'b0000000000000000;
       ph_real_24  <= 16'b0000000000000000;
       ph_real_25  <= 16'b0000000000000000;
       ph_real_26  <= 16'b0000000000000000;
       ph_real_27  <= 16'b0000000000000000;
       ph_real_28  <= 16'b0000000000000000;
       ph_real_29  <= 16'b0000000000000000;
       ph_real_30  <= 16'b0000000000000000;
       ph_real_31  <= 16'b0000000000000000;
       ph_real_32  <= 16'b0000000000000000;
       ph_real_33  <= 16'b0000000000000000;
       ph_real_34  <= 16'b0000000000000000;
       ph_real_35  <= 16'b0000000000000000; 
       ph_real_36  <= 16'b0000000000000000;
       ph_real_37  <= 16'b0000000000000000;
       ph_real_38  <= 16'b0000000000000000;
       ph_real_39  <= 16'b0000000000000000;
       ph_real_40  <= 16'b0000000000000000;
       ph_real_41  <= 16'b0000000000000000;
       ph_real_42  <= 16'b0000000000000000;
       ph_real_43  <= 16'b0000000000000000;
       ph_real_44  <= 16'b0000000000000000;
       ph_real_45  <= 16'b0000000000000000;
       ph_real_46  <= 16'b0000000000000000;
       ph_real_47  <= 16'b0000000000000000;
       ph_real_48  <= 16'b0000000000000000;
       
      ph_image_1 =  16'b0000000000000000;
      ph_image_2 =  16'b0000000000000000;
      ph_image_3 =  16'b0000000000000000; 
      ph_image_4 =  16'b0000000000000000;
      ph_image_5 =  16'b0000000000000000;
      ph_image_6 =  16'b0000000000000000;
      ph_image_7 =  16'b0000000000000000;
      ph_image_8 =  16'b0000000000000000;
      ph_image_9 =  16'b0000000000000000;
      ph_image_10<= 16'b0000000000000000;
      ph_image_11<= 16'b0000000000000000;
      ph_image_12<= 16'b0000000000000000;
      ph_image_13<= 16'b0000000000000000;
      ph_image_14<= 16'b0000000000000000;
      ph_image_15<= 16'b0000000000000000;
      ph_image_16<= 16'b0000000000000000;
      ph_image_17<= 16'b0000000000000000;
      ph_image_18<= 16'b0000000000000000;
      ph_image_19<= 16'b0000000000000000;
      ph_image_20<= 16'b0000000000000000;
      ph_image_21<= 16'b0000000000000000;
      ph_image_22<= 16'b0000000000000000;
      ph_image_23<= 16'b0000000000000000;
      ph_image_24<= 16'b0000000000000000;
      ph_image_25<= 16'b0000000000000000;
      ph_image_26<= 16'b0000000000000000;
      ph_image_27<= 16'b0000000000000000;
      ph_image_28<= 16'b0000000000000000;
      ph_image_29<= 16'b0000000000000000;
      ph_image_30<= 16'b0000000000000000;
      ph_image_31<= 16'b0000000000000000;
      ph_image_32<= 16'b0000000000000000;
      ph_image_33<= 16'b0000000000000000;
      ph_image_34<= 16'b0000000000000000;
      ph_image_35<= 16'b0000000000000000; 
      ph_image_36<= 16'b0000000000000000;
      ph_image_37<= 16'b0000000000000000;
      ph_image_38<= 16'b0000000000000000;
      ph_image_39<= 16'b0000000000000000;
      ph_image_40<= 16'b0000000000000000;
      ph_image_41<= 16'b0000000000000000;
      ph_image_42<= 16'b0000000000000000;
      ph_image_43<= 16'b0000000000000000;
      ph_image_44<= 16'b0000000000000000;
      ph_image_45<= 16'b0000000000000000;
      ph_image_46<= 16'b0000000000000000;
      ph_image_47<= 16'b0000000000000000;
      ph_image_48<= 16'b0000000000000000;
       end
    endcase
end





//dbf_phase_cormic dbf_phase_top_fangwei(
//    .clk(clk_120m),
    
//    .phase_data_1  (phase_data_1 ),
//    .phase_data_2  (phase_data_2 ),
//    .phase_data_3  (phase_data_3 ),
//    .phase_data_4  (phase_data_4 ),
//    .phase_data_5  (phase_data_5 ),
//    .phase_data_6  (phase_data_6 ),
//    .phase_data_7  (phase_data_7 ),
//    .phase_data_8  (phase_data_8 ),
//    .phase_data_9  (phase_data_9 ),
//    .phase_data_10 (phase_data_10 ),
//    .phase_data_11 (phase_data_11 ),
//    .phase_data_12 (phase_data_12 ),
//    .phase_data_13 (phase_data_13 ),
//    .phase_data_14 (phase_data_14 ),
//    .phase_data_15 (phase_data_15 ),
//    .phase_data_16 (phase_data_16 ),
//    .phase_data_17 (phase_data_17 ),
//    .phase_data_18 (phase_data_18 ),
//    .phase_data_19 (phase_data_19 ),
//    .phase_data_20 (phase_data_20 ),
//    .phase_data_21 (phase_data_21 ),
//    .phase_data_22 (phase_data_22 ),
//    .phase_data_23 (phase_data_23 ),
//    .phase_data_24 (phase_data_24 ),
//    .phase_data_25 (phase_data_25 ),
//    .phase_data_26 (phase_data_26 ),
//    .phase_data_27 (phase_data_27 ),
//    .phase_data_28 (phase_data_28 ),
//    .phase_data_29 (phase_data_29 ),
//    .phase_data_30 (phase_data_30 ),
//    .phase_data_31 (phase_data_31 ),
//    .phase_data_32 (phase_data_32 ),
//    .phase_data_33 (phase_data_33 ),
//    .phase_data_34 (phase_data_34 ),
//    .phase_data_35 (phase_data_35 ),
//    .phase_data_36 (phase_data_36 ),
//    .phase_data_37 (phase_data_37 ),
//    .phase_data_38 (phase_data_38 ),
//    .phase_data_39 (phase_data_39 ),
//    .phase_data_40 (phase_data_40 ),
//    .phase_data_41 (phase_data_41 ),
//    .phase_data_42 (phase_data_42 ),
//    .phase_data_43 (phase_data_43 ),
//    .phase_data_44 (phase_data_44 ),
//    .phase_data_45 (phase_data_45 ),
//    .phase_data_46 (phase_data_46 ),
//    .phase_data_47 (phase_data_47 ),
//    .phase_data_48 (phase_data_48 ),
   
    
//    .phase_data_valid(phase_data_valid),
    
    
//    .ph_real_1  (ph_real_1  ),
//    .ph_real_2  (ph_real_2  ),
//    .ph_real_3  (ph_real_3  ),
//    .ph_real_4  (ph_real_4  ),
//    .ph_real_5  (ph_real_5  ),
//    .ph_real_6  (ph_real_6  ),
//    .ph_real_7  (ph_real_7  ),
//    .ph_real_8  (ph_real_8  ),
//    .ph_real_9  (ph_real_9  ),
//    .ph_real_10 (ph_real_10 ),
//    .ph_real_11 (ph_real_11 ),
//    .ph_real_12 (ph_real_12 ),
//    .ph_real_13 (ph_real_13 ),
//    .ph_real_14 (ph_real_14 ),
//    .ph_real_15 (ph_real_15 ),
//    .ph_real_16 (ph_real_16 ),
//    .ph_real_17 (ph_real_17 ),
//    .ph_real_18 (ph_real_18 ),
//    .ph_real_19 (ph_real_19 ),
//    .ph_real_20 (ph_real_20 ),
//    .ph_real_21 (ph_real_21 ),
//    .ph_real_22 (ph_real_22 ),
//    .ph_real_23 (ph_real_23 ),
//    .ph_real_24 (ph_real_24 ),
//    .ph_real_25 (ph_real_25 ),
//    .ph_real_26 (ph_real_26 ),
//    .ph_real_27 (ph_real_27 ),
//    .ph_real_28 (ph_real_28 ),
//    .ph_real_29 (ph_real_29 ),
//    .ph_real_30 (ph_real_30 ),
//    .ph_real_31 (ph_real_31 ),
//    .ph_real_32 (ph_real_32 ),
//    .ph_real_33 (ph_real_33 ),
//    .ph_real_34 (ph_real_34 ),
//    .ph_real_35 (ph_real_35 ),
//    .ph_real_36 (ph_real_36 ),
//    .ph_real_37 (ph_real_37 ),
//    .ph_real_38 (ph_real_38 ),
//    .ph_real_39 (ph_real_39 ),
//    .ph_real_40 (ph_real_40 ),
//    .ph_real_41 (ph_real_41 ),
//    .ph_real_42 (ph_real_42 ),
//    .ph_real_43 (ph_real_43 ),
//    .ph_real_44 (ph_real_44 ),
//    .ph_real_45 (ph_real_45 ),
//    .ph_real_46 (ph_real_46 ),
//    .ph_real_47 (ph_real_47 ),
//    .ph_real_48 (ph_real_48 ),

    
    
//    .ph_image_1  (ph_image_1  ),
//    .ph_image_2  (ph_image_2  ),
//    .ph_image_3  (ph_image_3  ),
//    .ph_image_4  (ph_image_4  ),
//    .ph_image_5  (ph_image_5  ),
//    .ph_image_6  (ph_image_6  ),
//    .ph_image_7  (ph_image_7  ),
//    .ph_image_8  (ph_image_8  ),
//    .ph_image_9  (ph_image_9  ),
//    .ph_image_10 (ph_image_10 ),
//    .ph_image_11 (ph_image_11 ),
//    .ph_image_12 (ph_image_12 ),
//    .ph_image_13 (ph_image_13 ),
//    .ph_image_14 (ph_image_14 ),
//    .ph_image_15 (ph_image_15 ),
//    .ph_image_16 (ph_image_16 ),
//    .ph_image_17 (ph_image_17 ),
//    .ph_image_18 (ph_image_18 ),
//    .ph_image_19 (ph_image_19 ),
//    .ph_image_20 (ph_image_20 ),
//    .ph_image_21 (ph_image_21 ),
//    .ph_image_22 (ph_image_22 ),
//    .ph_image_23 (ph_image_23 ),
//    .ph_image_24 (ph_image_24 ),
//    .ph_image_25 (ph_image_25 ),
//    .ph_image_26 (ph_image_26 ),
//    .ph_image_27 (ph_image_27 ),
//    .ph_image_28 (ph_image_28 ),
//    .ph_image_29 (ph_image_29 ),
//    .ph_image_30 (ph_image_30 ),
//    .ph_image_31 (ph_image_31 ),
//    .ph_image_32 (ph_image_32 ),
//    .ph_image_33 (ph_image_33 ),
//    .ph_image_34 (ph_image_34 ),
//    .ph_image_35 (ph_image_35 ),
//    .ph_image_36 (ph_image_36 ),
//    .ph_image_37 (ph_image_37 ),
//    .ph_image_38 (ph_image_38 ),
//    .ph_image_39 (ph_image_39 ),
//    .ph_image_40 (ph_image_40 ),
//    .ph_image_41 (ph_image_41 ),
//    .ph_image_42 (ph_image_42 ),
//    .ph_image_43 (ph_image_43 ),
//    .ph_image_44 (ph_image_44 ),
//    .ph_image_45 (ph_image_45 ),
//    .ph_image_46 (ph_image_46 ),
//    .ph_image_47 (ph_image_47 ),
//    .ph_image_48 (ph_image_48 )

//    );
///////////////////////////////////////////////////////////////////////////
    wire [31:0]data_sum_I1; 
    wire [31:0]data_sum_Q1; 
    wire [31:0]data_sum_I2; 
    wire [31:0]data_sum_Q2; 
    wire [31:0]data_sum_I3; 
    wire [31:0]data_sum_Q3; 
    wire [31:0]data_sum_I4; 
    wire [31:0]data_sum_Q4; 
    wire [31:0]data_sum_I5; 
    wire [31:0]data_sum_Q5; 
    wire [31:0]data_sum_I6; 
    wire [31:0]data_sum_Q6; 
    wire [31:0]data_sum_I7; 
    wire [31:0]data_sum_Q7; 
    wire [31:0]data_sum_I8; 
    wire [31:0]data_sum_Q8; 
    wire [31:0]data_sum_I9; 
    wire [31:0]data_sum_Q9; 
    wire [31:0]data_sum_I10;
    wire [31:0]data_sum_Q10;
    wire [31:0]data_sum_I11;
    wire [31:0]data_sum_Q11;
    wire [31:0]data_sum_I12;
    wire [31:0]data_sum_Q12;
    wire [31:0]data_sum_I13;
    wire [31:0]data_sum_Q13;
    wire [31:0]data_sum_I14;
    wire [31:0]data_sum_Q14;
    wire [31:0]data_sum_I15;
    wire [31:0]data_sum_Q15;
    wire [31:0]data_sum_I16;
    wire [31:0]data_sum_Q16;
    wire [31:0]data_sum_I17; 
    wire [31:0]data_sum_Q17; 
    wire [31:0]data_sum_I18;
    wire [31:0]data_sum_Q18;
    wire [31:0]data_sum_I19;
    wire [31:0]data_sum_Q19;
    wire [31:0]data_sum_I20;
    wire [31:0]data_sum_Q20;
    wire [31:0]data_sum_I21;
    wire [31:0]data_sum_Q21;
    wire [31:0]data_sum_I22;
    wire [31:0]data_sum_Q22;
    wire [31:0]data_sum_I23;
    wire [31:0]data_sum_Q23;
    wire [31:0]data_sum_I24;
    wire [31:0]data_sum_Q24;


dbf_v1 add_1_24(
        .clk(clk_120m),
        .dataI(dataI),
        .dataQ(dataQ),
        .data_in_valid(data_in_valid),
        .fw_cut_ctl(fw_cut_ctl),
        
    .ph_real_1  (ph_real_1  ),
    .ph_real_2  (ph_real_2  ),
    .ph_real_3  (ph_real_3  ),
    .ph_real_4  (ph_real_4  ),
    .ph_real_5  (ph_real_5  ),
    .ph_real_6  (ph_real_6  ),
    .ph_real_7  (ph_real_7  ),
    .ph_real_8  (ph_real_8  ),
    .ph_real_9  (ph_real_9  ),
    .ph_real_10 (ph_real_10 ),
    .ph_real_11 (ph_real_11 ),
    .ph_real_12 (ph_real_12 ),
    .ph_real_13 (ph_real_13 ),
    .ph_real_14 (ph_real_14 ),
    .ph_real_15 (ph_real_15 ),
    .ph_real_16 (ph_real_16 ),
    .ph_real_17 (ph_real_17 ),
    .ph_real_18 (ph_real_18 ),
    .ph_real_19 (ph_real_19 ),
    .ph_real_20 (ph_real_20 ),
    .ph_real_21 (ph_real_21 ),
    .ph_real_22 (ph_real_22 ),
    .ph_real_23 (ph_real_23 ),
    .ph_real_24 (ph_real_24 ),
    .ph_image_1  (ph_image_1  ),
    .ph_image_2  (ph_image_2  ),
    .ph_image_3  (ph_image_3  ),
    .ph_image_4  (ph_image_4  ),
    .ph_image_5  (ph_image_5  ),
    .ph_image_6  (ph_image_6  ),
    .ph_image_7  (ph_image_7  ),
    .ph_image_8  (ph_image_8  ),
    .ph_image_9  (ph_image_9  ),
    .ph_image_10 (ph_image_10 ),
    .ph_image_11 (ph_image_11 ),
    .ph_image_12 (ph_image_12 ),
    .ph_image_13 (ph_image_13 ),
    .ph_image_14 (ph_image_14 ),
    .ph_image_15 (ph_image_15 ),
    .ph_image_16 (ph_image_16 ),
    .ph_image_17 (ph_image_17 ),
    .ph_image_18 (ph_image_18 ),
    .ph_image_19 (ph_image_19 ),
    .ph_image_20 (ph_image_20 ),
    .ph_image_21 (ph_image_21 ),
    .ph_image_22 (ph_image_22 ),
    .ph_image_23 (ph_image_23 ),
    .ph_image_24 (ph_image_24 ),
    
        .A_1 (A_1 ),
        .A_2 (A_2 ),
        .A_3 (A_3 ),
        .A_4 (A_4 ),
        .A_5 (A_5 ),
        .A_6 (A_6 ),
        .A_7 (A_7 ),
        .A_8 (A_8 ),
        .A_9 (A_9 ),
        .A_10(A_10),
        .A_11(A_11),
        .A_12(A_12),
        .A_13(A_13),
        .A_14(A_14),
        .A_15(A_15),
        .A_16(A_16),
        .A_17(A_17),
        .A_18(A_18),
        .A_19(A_19),
        .A_20(A_20),
        .A_21(A_21),
        .A_22(A_22),
        .A_23(A_23),
        .A_24(A_24),
        
       
        
        .phase_data_valid(phase_data_valid),
        
        .add_out_I(add_out_1_24_I),
        .add_out_Q(add_out_1_24_Q),
        .data_out_valid_1(data_out_valid),
        
        .data_sum_I1(data_sum_I1),
        .data_sum_Q1(data_sum_Q1),
        .data_sum_I2(data_sum_I2),
        .data_sum_Q2(data_sum_Q2),
        .data_sum_I3(data_sum_I3),
        .data_sum_Q3(data_sum_Q3),
        .data_sum_I4(data_sum_I4),
        .data_sum_Q4(data_sum_Q4),
        .data_sum_I5(data_sum_I5),
        .data_sum_Q5(data_sum_Q5),
        .data_sum_I6(data_sum_I6),
        .data_sum_Q6(data_sum_Q6),
        .data_sum_I7(data_sum_I7),
        .data_sum_Q7(data_sum_Q7),
        .data_sum_I8(data_sum_I8),
        .data_sum_Q8(data_sum_Q8),
        .data_sum_I9(data_sum_I9),
        .data_sum_Q9(data_sum_Q9),
        .data_sum_I10(data_sum_I10),
        .data_sum_Q10(data_sum_Q10),
        .data_sum_I11(data_sum_I11),
        .data_sum_Q11(data_sum_Q11),
        .data_sum_I12(data_sum_I12),
        .data_sum_Q12(data_sum_Q12),
        .data_sum_I13(data_sum_I13),
        .data_sum_Q13(data_sum_Q13),
        .data_sum_I14(data_sum_I14),
        .data_sum_Q14(data_sum_Q14),
        .data_sum_I15(data_sum_I15),
        .data_sum_Q15(data_sum_Q15),
        .data_sum_I16(data_sum_I16),
        .data_sum_Q16(data_sum_Q16),
        .data_sum_I17(data_sum_I17),
        .data_sum_Q17(data_sum_Q17),
        .data_sum_I18(data_sum_I18),
        .data_sum_Q18(data_sum_Q18),
        .data_sum_I19(data_sum_I19),
        .data_sum_Q19(data_sum_Q19),
        .data_sum_I20(data_sum_I20),
        .data_sum_Q20(data_sum_Q20),
        .data_sum_I21(data_sum_I21),
        .data_sum_Q21(data_sum_Q21),
        .data_sum_I22(data_sum_I22),
        .data_sum_Q22(data_sum_Q22),
        .data_sum_I23(data_sum_I23),
        .data_sum_Q23(data_sum_Q23),
        .data_sum_I24(data_sum_I24),
        .data_sum_Q24(data_sum_Q24)     
  
);


wire [31:0]data_sum_I25;
wire [31:0]data_sum_Q25;
wire [31:0]data_sum_I26;
wire [31:0]data_sum_Q26;
wire [31:0]data_sum_I27;
wire [31:0]data_sum_Q27;
wire [31:0]data_sum_I28;
wire [31:0]data_sum_Q28;
wire [31:0]data_sum_I29;
wire [31:0]data_sum_Q29;
wire [31:0]data_sum_I30;
wire [31:0]data_sum_Q30;
wire [31:0]data_sum_I31;
wire [31:0]data_sum_Q31;
wire [31:0]data_sum_I32;
wire [31:0]data_sum_Q32;
wire [31:0]data_sum_I33;
wire [31:0]data_sum_Q33;
wire [31:0]data_sum_I34;
wire [31:0]data_sum_Q34;
wire [31:0]data_sum_I35;
wire [31:0]data_sum_Q35;
wire [31:0]data_sum_I36;
wire [31:0]data_sum_Q36;
wire [31:0]data_sum_I37;
wire [31:0]data_sum_Q37;
wire [31:0]data_sum_I38;
wire [31:0]data_sum_Q38;
wire [31:0]data_sum_I39;
wire [31:0]data_sum_Q39;
wire [31:0]data_sum_I40;
wire [31:0]data_sum_Q40;
wire [31:0]data_sum_I41;
wire [31:0]data_sum_Q41;
wire [31:0]data_sum_I42;
wire [31:0]data_sum_Q42;
wire [31:0]data_sum_I43;
wire [31:0]data_sum_Q43;
wire [31:0]data_sum_I44;
wire [31:0]data_sum_Q44;
wire [31:0]data_sum_I45;
wire [31:0]data_sum_Q45;
wire [31:0]data_sum_I46;
wire [31:0]data_sum_Q46;
wire [31:0]data_sum_I47;
wire [31:0]data_sum_Q47;
wire [31:0]data_sum_I48;
wire [31:0]data_sum_Q48;


dbf_v1 add_25_48(
        .clk(clk_120m),
        .dataI(dataI),
        .dataQ(dataQ),
        .data_in_valid(data_in_valid),
        .fw_cut_ctl(fw_cut_ctl),
        
    .ph_real_1   (ph_real_25 ),
    .ph_real_2   (ph_real_26 ),
    .ph_real_3   (ph_real_27 ),
    .ph_real_4   (ph_real_28 ),
    .ph_real_5   (ph_real_29 ),
    .ph_real_6   (ph_real_30 ),
    .ph_real_7   (ph_real_31 ),
    .ph_real_8   (ph_real_32 ),
    .ph_real_9   (ph_real_33 ),
    .ph_real_10  (ph_real_34 ),
    .ph_real_11  (ph_real_35 ),
    .ph_real_12  (ph_real_36 ),
    .ph_real_13  (ph_real_37 ),
    .ph_real_14  (ph_real_38 ),
    .ph_real_15  (ph_real_39 ),
    .ph_real_16  (ph_real_40 ),
    .ph_real_17  (ph_real_41 ),
    .ph_real_18  (ph_real_42 ),
    .ph_real_19  (ph_real_43 ),
    .ph_real_20  (ph_real_44 ),
    .ph_real_21  (ph_real_45 ),
    .ph_real_22  (ph_real_46 ),
    .ph_real_23  (ph_real_47 ),
    .ph_real_24  (ph_real_48 ),
    .ph_image_1  (ph_image_25 ),
    .ph_image_2  (ph_image_26 ),
    .ph_image_3  (ph_image_27 ),
    .ph_image_4  (ph_image_28 ),
    .ph_image_5  (ph_image_29 ),
    .ph_image_6  (ph_image_30 ),
    .ph_image_7  (ph_image_31 ),
    .ph_image_8  (ph_image_32 ),
    .ph_image_9  (ph_image_33 ),
    .ph_image_10 (ph_image_34 ),
    .ph_image_11 (ph_image_35 ),
    .ph_image_12 (ph_image_36 ),
    .ph_image_13 (ph_image_37 ),
    .ph_image_14 (ph_image_38 ),
    .ph_image_15 (ph_image_39 ),
    .ph_image_16 (ph_image_40 ),
    .ph_image_17 (ph_image_41 ),
    .ph_image_18 (ph_image_42 ),
    .ph_image_19 (ph_image_43 ),
    .ph_image_20 (ph_image_44 ),
    .ph_image_21 (ph_image_45 ),
    .ph_image_22 (ph_image_46 ),
    .ph_image_23 (ph_image_47 ),
    .ph_image_24 (ph_image_48 ),
    
        .A_1 (A_25),
        .A_2 (A_26),
        .A_3 (A_27),
        .A_4 (A_28),
        .A_5 (A_29),
        .A_6 (A_30),
        .A_7 (A_31),
        .A_8 (A_32),
        .A_9 (A_33),
        .A_10(A_34),
        .A_11(A_35),
        .A_12(A_36),
        .A_13(A_37),
        .A_14(A_38),
        .A_15(A_39),
        .A_16(A_40),
        .A_17(A_41),
        .A_18(A_42),
        .A_19(A_43),
        .A_20(A_44),
        .A_21(A_45),
        .A_22(A_46),
        .A_23(A_47),
        .A_24(A_48),

        
       
        .phase_data_valid(phase_data_valid),
        
        .add_out_I(add_out_25_48_I),
        .add_out_Q(add_out_25_48_Q),
        .data_out_valid_1(),
        
        .data_sum_I1(data_sum_I25),
        .data_sum_Q1(data_sum_Q25),
        .data_sum_I2(data_sum_I26),
        .data_sum_Q2(data_sum_Q26),
        .data_sum_I3(data_sum_I27),
        .data_sum_Q3(data_sum_Q27),
        .data_sum_I4(data_sum_I28),
        .data_sum_Q4(data_sum_Q28),
        .data_sum_I5(data_sum_I29),
        .data_sum_Q5(data_sum_Q29),
        .data_sum_I6(data_sum_I30),
        .data_sum_Q6(data_sum_Q30),
        .data_sum_I7(data_sum_I31),
        .data_sum_Q7(data_sum_Q31),
        .data_sum_I8(data_sum_I32),
        .data_sum_Q8(data_sum_Q32),
        .data_sum_I9(data_sum_I33),
        .data_sum_Q9(data_sum_Q33),
        .data_sum_I10(data_sum_I34),
        .data_sum_Q10(data_sum_Q34),
        .data_sum_I11(data_sum_I35),
        .data_sum_Q11(data_sum_Q35),
        .data_sum_I12(data_sum_I36),
        .data_sum_Q12(data_sum_Q36),
        .data_sum_I13(data_sum_I37),
        .data_sum_Q13(data_sum_Q37),
        .data_sum_I14(data_sum_I38),
        .data_sum_Q14(data_sum_Q38),
        .data_sum_I15(data_sum_I39),
        .data_sum_Q15(data_sum_Q39),
        .data_sum_I16(data_sum_I40),
        .data_sum_Q16(data_sum_Q40),
        .data_sum_I17(data_sum_I41),   
        .data_sum_Q17(data_sum_Q41),
        .data_sum_I18(data_sum_I42),
        .data_sum_Q18(data_sum_Q42),
        .data_sum_I19(data_sum_I43),
        .data_sum_Q19(data_sum_Q43),
        .data_sum_I20(data_sum_I44),
        .data_sum_Q20(data_sum_Q44),
        .data_sum_I21(data_sum_I45),
        .data_sum_Q21(data_sum_Q45),
        .data_sum_I22(data_sum_I46),
        .data_sum_Q22(data_sum_Q46),
        .data_sum_I23(data_sum_I47),
        .data_sum_Q23(data_sum_Q47),
        .data_sum_I24(data_sum_I48),
        .data_sum_Q24(data_sum_Q48)
       
          
);
    
//ila_fangweisub ila_fangweisub_1 (
//	.clk(clk_120m), // input wire clk


//	.probe0 (data_sum_I1), // input wire [31:0]  probe0  
//	.probe1 (data_sum_Q1), // input wire [31:0]  probe1 
//	.probe2 (data_sum_I2), // input wire [31:0]  probe2 
//	.probe3 (data_sum_Q2), // input wire [31:0]  probe3 
//	.probe4 (data_sum_I3), // input wire [31:0]  probe4 
//	.probe5 (data_sum_Q3), // input wire [31:0]  probe5 
//	.probe6 (data_sum_I4), // input wire [31:0]  probe6 
//	.probe7 (data_sum_Q4), // input wire [31:0]  probe7 
//	.probe8 (data_sum_I5), // input wire [31:0]  probe8 
//	.probe9 (data_sum_Q5), // input wire [31:0]  probe9 
//	.probe10(data_sum_I6), // input wire [31:0]  probe10 
//	.probe11(data_sum_Q6), // input wire [31:0]  probe11 
//	.probe12(data_sum_I7), // input wire [31:0]  probe12 
//	.probe13(data_sum_Q7), // input wire [31:0]  probe13 
//	.probe14(data_sum_I8), // input wire [31:0]  probe14 
//	.probe15(data_sum_Q8), // input wire [31:0]  probe15 
//	.probe16(data_sum_I9), // input wire [31:0]  probe16 
//	.probe17(data_sum_Q9), // input wire [31:0]  probe17 
//	.probe18(data_sum_I10), // input wire [31:0]  probe18 
//	.probe19(data_sum_Q10), // input wire [31:0]  probe19 
//	.probe20(data_sum_I11), // input wire [31:0]  probe20 
//	.probe21(data_sum_Q11), // input wire [31:0]  probe21 
//	.probe22(data_sum_I12), // input wire [31:0]  probe22 
//	.probe23(data_sum_Q12), // input wire [31:0]  probe23 
//	.probe24(data_sum_I13), // input wire [31:0]  probe24 
//	.probe25(data_sum_Q13), // input wire [31:0]  probe25 
//	.probe26(data_sum_I14), // input wire [31:0]  probe26 
//	.probe27(data_sum_Q14), // input wire [31:0]  probe27 
//	.probe28(data_sum_I15), // input wire [31:0]  probe28 
//	.probe29(data_sum_Q15), // input wire [31:0]  probe29 
//	.probe30(data_sum_I16), // input wire [31:0]  probe30 
//	.probe31(data_sum_Q16), // input wire [31:0]  probe31 
//	.probe32(data_sum_I17), // input wire [31:0]  probe32 
//	.probe33(data_sum_Q17), // input wire [31:0]  probe33 
//	.probe34(data_sum_I18), // input wire [31:0]  probe34 
//	.probe35(data_sum_Q18), // input wire [31:0]  probe35 
//	.probe36(data_sum_I19), // input wire [31:0]  probe36 
//	.probe37(data_sum_Q19), // input wire [31:0]  probe37 
//	.probe38(data_sum_I20), // input wire [31:0]  probe38 
//	.probe39(data_sum_Q20), // input wire [31:0]  probe39 
//	.probe40(data_sum_I21), // input wire [31:0]  probe40 
//	.probe41(data_sum_Q21), // input wire [31:0]  probe41 
//	.probe42(data_sum_I22), // input wire [31:0]  probe42 
//	.probe43(data_sum_Q22), // input wire [31:0]  probe43 
//	.probe44(data_sum_I23), // input wire [31:0]  probe44 
//	.probe45(data_sum_Q23), // input wire [31:0]  probe45 
//	.probe46(data_sum_I24), // input wire [31:0]  probe46 
//	.probe47(data_sum_Q24), // input wire [31:0]  probe47 
//	.probe48(data_sum_I25), // input wire [31:0]  probe48 
//	.probe49(data_sum_Q25), // input wire [31:0]  probe49 
//	.probe50(data_sum_I26), // input wire [31:0]  probe50 
//	.probe51(data_sum_Q26), // input wire [31:0]  probe51 
//	.probe52(data_sum_I27), // input wire [31:0]  probe52 
//	.probe53(data_sum_Q27), // input wire [31:0]  probe53 
//	.probe54(data_sum_I28), // input wire [31:0]  probe54 
//	.probe55(data_sum_Q28), // input wire [31:0]  probe55 
//	.probe56(data_sum_I29), // input wire [31:0]  probe56 
//	.probe57(data_sum_Q29), // input wire [31:0]  probe57 
//	.probe58(data_sum_I30), // input wire [31:0]  probe58 
//	.probe59(data_sum_Q30), // input wire [31:0]  probe59 
//	.probe60(data_sum_I31), // input wire [31:0]  probe60 
//	.probe61(data_sum_Q31), // input wire [31:0]  probe61 
//	.probe62(data_sum_I32), // input wire [31:0]  probe62 
//	.probe63(data_sum_Q32) // input wire [31:0]  probe63
	
//);


//ila_4 fw_t (
//	.clk(clk_120m), // input wire clk

//	.probe0(dataI), // input wire [15:0]  probe0  
//	.probe1(dataQ), // input wire [15:0]  probe1 
//	.probe2(data_in_valid), // input wire [0:0]  probe2 
//	.probe3(fpga_gpio), // input wire [15:0]  probe3 
//	.probe4(add_out_1_24_I), // input wire [15:0]  probe4 
//	.probe5(add_out_1_24_Q), // input wire [15:0]  probe5 
//	.probe6(add_out_25_48_I), // input wire [15:0]  probe6 
//	.probe7(add_out_25_48_Q), // input wire [15:0]  probe7 
//	.probe8(data_out_valid) // input wire [0:0]  probe8 
	
	
	
	
//);

//ila_2 FW_PH (
//	.clk(clk_120m), // input wire clk


//	.probe0(phase_data_1), // input wire [15:0]  probe0  
//	.probe1(phase_data_2), // input wire [15:0]  probe1 
//	.probe2(phase_data_3), // input wire [15:0]  probe2 
//	.probe3(phase_data_4), // input wire [15:0]  probe3 
//	.probe4(phase_data_5), // input wire [15:0]  probe4 
//	.probe5(phase_data_6), // input wire [15:0]  probe5 
//	.probe6(phase_data_7), // input wire [15:0]  probe6 
//	.probe7(phase_data_8), // input wire [15:0]  probe7 
//	.probe8(phase_data_9), // input wire [15:0]  probe8 
//	.probe9(phase_data_10), // input wire [15:0]  probe9 
//	.probe10(phase_data_11), // input wire [15:0]  probe10 
//	.probe11(phase_data_12), // input wire [15:0]  probe11 
//	.probe12(phase_data_13), // input wire [15:0]  probe12 
//	.probe13(phase_data_14), // input wire [15:0]  probe13 
//	.probe14(phase_data_15), // input wire [15:0]  probe14 
//	.probe15(phase_data_16), // input wire [15:0]  probe15 
//	.probe16(phase_data_17), // input wire [15:0]  probe16 
//	.probe17(phase_data_18), // input wire [15:0]  probe17 
//	.probe18(phase_data_19), // input wire [15:0]  probe18 
//	.probe19(phase_data_20), // input wire [15:0]  probe19 
//	.probe20(phase_data_21), // input wire [15:0]  probe20 
//	.probe21(phase_data_22), // input wire [15:0]  probe21 
//	.probe22(phase_data_23), // input wire [15:0]  probe22 
//	.probe23(phase_data_24), // input wire [15:0]  probe23 
//	.probe24(phase_data_25), // input wire [15:0]  probe24 
//	.probe25(phase_data_26), // input wire [15:0]  probe25 
//	.probe26(phase_data_27), // input wire [15:0]  probe26 
//	.probe27(phase_data_28), // input wire [15:0]  probe27 
//	.probe28(phase_data_29), // input wire [15:0]  probe28 
//	.probe29(phase_data_30), // input wire [15:0]  probe29 
//	.probe30(phase_data_31), // input wire [15:0]  probe30 
//	.probe31(phase_data_32) // input wire [15:0]  probe31
//);           
//ila_pd_fangwei ila_pd_fangwei_1 (
//	.clk(clk_120m), // input wire clk


//	.probe0(ph_real_1), // input wire [15:0]  probe0  
//	.probe1(ph_real_2), // input wire [15:0]  probe1 
//	.probe2(ph_real_3), // input wire [15:0]  probe2 
//	.probe3(ph_real_4), // input wire [15:0]  probe3 
//	.probe4(ph_real_5), // input wire [15:0]  probe4 
//	.probe5(ph_real_6), // input wire [15:0]  probe5 
//	.probe6(ph_real_7), // input wire [15:0]  probe6 
//	.probe7(ph_real_8), // input wire [15:0]  probe7 
//	.probe8(ph_real_9), // input wire [15:0]  probe8 
//	.probe9(ph_real_10), // input wire [15:0]  probe9 
//	.probe10(ph_real_11), // input wire [15:0]  probe10 
//	.probe11(ph_real_12), // input wire [15:0]  probe11 
//	.probe12(ph_real_13), // input wire [15:0]  probe12 
//	.probe13(ph_real_14), // input wire [15:0]  probe13 
//	.probe14(ph_real_15), // input wire [15:0]  probe14 
//	.probe15(ph_real_16), // input wire [15:0]  probe15 
//	.probe16(ph_real_17), // input wire [15:0]  probe16 
//	.probe17(ph_real_18), // input wire [15:0]  probe17 
//	.probe18(ph_real_19), // input wire [15:0]  probe18 
//	.probe19(ph_real_20), // input wire [15:0]  probe19 
//	.probe20(ph_real_21), // input wire [15:0]  probe20 
//	.probe21(ph_real_22), // input wire [15:0]  probe21 
//	.probe22(ph_real_23), // input wire [15:0]  probe22 
//	.probe23(ph_real_24), // input wire [15:0]  probe23 
//	.probe24(ph_real_25), // input wire [15:0]  probe24 
//	.probe25(ph_real_26), // input wire [15:0]  probe25 
//	.probe26(ph_real_27), // input wire [15:0]  probe26 
//	.probe27(ph_real_28), // input wire [15:0]  probe27 
//	.probe28(ph_real_29), // input wire [15:0]  probe28 
//	.probe29(ph_real_30), // input wire [15:0]  probe29 
//	.probe30(ph_real_31), // input wire [15:0]  probe30 
//	.probe31(ph_real_32), // input wire [15:0]  probe31 
//	.probe32(ph_real_33), // input wire [15:0]  probe32 
//	.probe33(ph_real_34), // input wire [15:0]  probe33 
//	.probe34(ph_real_35), // input wire [15:0]  probe34 
//	.probe35(ph_real_36), // input wire [15:0]  probe35 
//	.probe36(ph_real_37), // input wire [15:0]  probe36 
//	.probe37(ph_real_38), // input wire [15:0]  probe37 
//	.probe38(ph_real_39), // input wire [15:0]  probe38 
//	.probe39(ph_real_40), // input wire [15:0]  probe39 
//	.probe40(ph_real_41), // input wire [15:0]  probe40 
//	.probe41(ph_real_42), // input wire [15:0]  probe41 
//	.probe42(ph_real_43), // input wire [15:0]  probe42 
//	.probe43(ph_real_44), // input wire [15:0]  probe43 
//	.probe44(ph_real_45), // input wire [15:0]  probe44 
//	.probe45(ph_real_46), // input wire [15:0]  probe45 
//	.probe46(ph_real_47), // input wire [15:0]  probe46 
//	.probe47(ph_real_48) // input wire [15:0]  probe47
//);
////ila_pd_fangwei ila_pd_fangwei_2 (
////	.clk(clk_120m), // input wire clk


//	.probe0(ph_image_1), // input wire [15:0]  probe0  
//	.probe1(ph_image_2), // input wire [15:0]  probe1 
//	.probe2(ph_image_3), // input wire [15:0]  probe2 
//	.probe3(ph_image_4), // input wire [15:0]  probe3 
//	.probe4(ph_image_5), // input wire [15:0]  probe4 
//	.probe5(ph_image_6), // input wire [15:0]  probe5 
//	.probe6(ph_image_7), // input wire [15:0]  probe6 
//	.probe7(ph_image_8), // input wire [15:0]  probe7 
//	.probe8(ph_image_9), // input wire [15:0]  probe8 
//	.probe9(ph_image_10), // input wire [15:0]  probe9 
//	.probe10(ph_image_11), // input wire [15:0]  probe10 
//	.probe11(ph_image_12), // input wire [15:0]  probe11 
//	.probe12(ph_image_13), // input wire [15:0]  probe12 
//	.probe13(ph_image_14), // input wire [15:0]  probe13 
//	.probe14(ph_image_15), // input wire [15:0]  probe14 
//	.probe15(ph_image_16), // input wire [15:0]  probe15 
//	.probe16(ph_image_17), // input wire [15:0]  probe16 
//	.probe17(ph_image_18), // input wire [15:0]  probe17 
//	.probe18(ph_image_19), // input wire [15:0]  probe18 
//	.probe19(ph_image_20), // input wire [15:0]  probe19 
//	.probe20(ph_image_21), // input wire [15:0]  probe20 
//	.probe21(ph_image_22), // input wire [15:0]  probe21 
//	.probe22(ph_image_23), // input wire [15:0]  probe22 
//	.probe23(ph_image_24), // input wire [15:0]  probe23 
//	.probe24(ph_image_25), // input wire [15:0]  probe24 
//	.probe25(ph_image_26), // input wire [15:0]  probe25 
//	.probe26(ph_image_27), // input wire [15:0]  probe26 
//	.probe27(ph_image_28), // input wire [15:0]  probe27 
//	.probe28(ph_image_29), // input wire [15:0]  probe28 
//	.probe29(ph_image_30), // input wire [15:0]  probe29 
//	.probe30(ph_image_31), // input wire [15:0]  probe30 
//	.probe31(ph_image_32), // input wire [15:0]  probe31 
//	.probe32(ph_image_33), // input wire [15:0]  probe32 
//	.probe33(ph_image_34), // input wire [15:0]  probe33 
//	.probe34(ph_image_35), // input wire [15:0]  probe34 
//	.probe35(ph_image_36), // input wire [15:0]  probe35 
//	.probe36(ph_image_37), // input wire [15:0]  probe36 
//	.probe37(ph_image_38), // input wire [15:0]  probe37 
//	.probe38(ph_image_39), // input wire [15:0]  probe38 
//	.probe39(ph_image_40), // input wire [15:0]  probe39 
//	.probe40(ph_image_41), // input wire [15:0]  probe40 
//	.probe41(ph_image_42), // input wire [15:0]  probe41 
//	.probe42(ph_image_43), // input wire [15:0]  probe42 
//	.probe43(ph_image_44), // input wire [15:0]  probe43 
//	.probe44(ph_image_45), // input wire [15:0]  probe44 
//	.probe45(ph_image_46), // input wire [15:0]  probe45 
//	.probe46(ph_image_47), // input wire [15:0]  probe46 
//	.probe47(ph_image_48) // input wire [15:0]  probe47
//);
    
endmodule
